��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P����z��{}H���_Q�hФ���]xy�0�|s��9߼L���حe=�3�����Uh=8G%�t���n�4��D�cm��zۜq�a��?w}HC�#u¨�`�L�Cަg
WS�1f�k��Z�W�Ԕa� �����O:_�ڋ"���Pܣ=2UܪWݒ%��u���!����?`Ӥ��T��(i'��}t�	Zje��tF��AB�.��v�4�`��U���� ۑ�梎n&�Y�m"�M a������W1ԍ��;&GM��=,	(�x��E�d�E��v�p������`v�Sn��%�p?��!��8�a���)1���Τ�L���6��.�� �(jO6��A)t(K� oR���)���P�h��a5M��V�N����Q6F<~���^ò��"�ic�0���.���{��1���kl��ߛ;��_��|�=�Uޅ�q�=�Ψ�	r��q
����_���,ͦ���z?�bj!x�Ǐ�<�+e�9���P]�CM�����åcY���J]�w6��9$���e�f~*�hk���~5W�f�E����RT����Ϗ4�RN>�1��_��(�{���.,��R�P:���X�/�W�!�C�S��X�F�� R?����h<?�Y�aPһ����'@M��s��9��e^�¨f�x
#p���&�N+ [�nL��*�һ�Hd���Hl���H��A��i�⃋��O!�Q����%�C�8�hz���]�˷	�n`�T�\��D
��j�2��qZ�P'�fk�W��&
���?�Y��� u���)�hڿ�����N�l�&P�h�P�Lg�?I^�Ob.Qܵ������w���ѫ�/s7r�=����"xX�zN,8���<�,8s	���A�b�5�o�@��b%k�br𲊐i���Y�6P����Tk!u�i�����+j]P��EF�(-��vz�4æl3�n1� ��I@��f�q��ɞh ����S�9;���v"�z�
�`c2r�ο5_�6��_
��i,�v
��,�����J�Y�<C�67YUZR�"y�W1�/Q`R�l�
0`�.sW�&L�ɷ�f��
�� ���Qh�@��k�v;�y�T*GLI=?d�B�B&- �lYP���Y�&�rP>�A[�Ş�cެ���\�Pc��T§{�<�v�M"8��	NI�H���9Ґ `	c�?\�����6�8}g֞�vҧ�|(��6�ǜ{H^�a�9Bl��8ܲ��q-Y�tld�z����j�Uh�և���l��e䅅�6��>Rk�U��9����d�<^�?`S��.?Z���o�ę3��52��>�bBeI�Q �󧒝ۧ�-�n5�e��?�j�{��@�*�X�h�0�e�����+��7�dr��d8j�^�����M�[50����o��V�lB���5�(�ڇp�O�U=��)f�N'������>:y
:״d��Q�ާ�&�0�#o~��&��O��S��Υ��րx�z}��4�^0��q�~L��I� ���bԜ�j�<-z�}��j=5v#9f�_|z��/M��X��ƀ�����c�3�̪�[���������m�� ~�� w��J� ^���"��2h��c
n�����#�`��/0��$l!�5ֈ":)�|����]
�R�@kB��?�ZN<�*���Ff��J�'�pS]`�Q��O�C��/A�>ړ�x�A�s$����\�]����>�PƱE�u٨��}�����n�JRݭ�=t��ېb�d�ǙP%�)W��x��6�cQ���O���aR�!�b?^l�ZQJ�1C����`ʽ��<a�+�O����@�g}�S�oR�3��*����z��SO���
�۽6#!�ۅC{Qoި�sAp�i�Ncʭ��m�T���L��C7��\��uD ��H�8��/��������KH~�f