��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd����a�n��>�ԍ�O�xjt���>�Qm�<�v`�������/�)�=���0A iʵ��	z+Lк�����vuk��vz��@I3j�����m�z#��-$z��uA�So����������0C�J�t�m��%գTF�����y�ǧ���wu����;�s�U�k���/{��	x,���@a�W4U���l��qL��
ki�PMf����ǐK�	���A�f�-߻v�ޑ����񿞜n��|�<m�LB,n�	Q�xA1 R��'�p�T-oYBV�4�=V�z��l���T��f�H):�'�r��XZA��	�(:*��Z�c+?��\O ��O{jC��[��İ�D�N}&s!��RK���ے�2Ƃ� �o�Z�5j@�pq�=����VX���#���;4����z diDm�k>P��A
�Hj��@����ޖè<�r8�r��ZZ4���DΪ��B�,H��:;8â�]:(�Dk��)s�E�%Kt��dL��A��R��"<�Y�󞠝�{A�~s�F~YYTn����*���G^�J?�鍒R��]o$!&���{2)�_���<I7���B�3/�eU�R"��;p��G��n�r$�Y�2�zz@��ST��)�&4�z�^�cs�I��`  4S�s�3*��
+��B��W
�s&Y��,�q$3HRs	Y��X��,��'я��T=���%  z���{J��8��l�����rNԙ��3���M2ºQ9~b�HD���ubկ["3TġD?Eylh����Hs�f��o�8=�J
�^�]|u�2���=_���������.��x��t;�n��9��N5���V��u�$C���G�͛��:�"8Þ_/ƄZ_�f�h�%:����ʵo��v�6o`��q�� h$�^����^�+����s���l���	j��1�l�P����N(鴄�9�� �h6�/V�Nӕ\�Hx�l�p�0l$q��G�7B�!������[O��\B3��K�-�Yu�J��/�������^S�]�A�+�EkBy��X(I�O�BE����%~rk�>����X���Dz%o]�H�s1��[����\�NR&�G0��w'D)N@�r�#S�`�>.E�[���ڱ�g�V�N��S���ݫ�����'�d�z����ψ\-����@��{)��)�����!;#�&�]�ڠ�>V���X��<������S]�^B��2���i50#�0z
��r�0�jm��x��$�lEo$�:�j��qc�@��B,$�D���n|8;k�#+{��}f��:E��\�i�@#��AC&���Z�7����s�8��9FPw����_�#�ܟo��{�=�E6��Q�]j�X=��V#�+�i �*��R���|�f�*+�"$��4`��o,����ˏ�	ʴ�̛��)�R��܃ذ*;̭¢����;b�ihQ��nF����<H:4�|�?�����{4� ���8|��}�ϡU濵9z�� ;�Z�+��ђH��`�J:�N�@�o�G����J��x��ҥ�*p�~�}��-�pc>�n����TJ˗FSE	�G<�K�Fc���+����81oR�,��T�9 �n(���VEP'g^�S}��B!�'L���fM���8
��j�p�A`u���V��k [�%�X���7Ր{��vp��o\��ud ��;��f��`)�H�d��-9�$3���[�t7��q�*������/��z�H~��M�܉�ߏ�zMt�φ^�Y�G�Sl���c6�"V���ǡ�3�d=�-����-�+�����`P����v�o����ĩ*tTR<��ח��ݮA{��}����$�;=���X��o}����A��d��;����T��aG���V�!� $͸)-)Tץ�.���:��y���9abPwe*�	ȦF\\��|���V��79ǉ����H")ޒCkYK�[RWD&�_Gn��D�&���pXXC	Ē���?d�ӧ���`�'��V8�l�TW�.rtr?\�\D����jk$����;`y�Іs� �����?�t�"B��9�T<Isuw�X`�	�XD���e�p�%��~�u��I����::�m
NߚT�W��]�Z���m�2��.��`�!��Y�����&�:���3>a��pB��@��,T�x!���{��(��(�EE���b����$`���g��q�Юp�������0�����N�9�m�4��J�4�����"��I-&z�y86 O�k�J[XdbC#;���1F�^-eդ��f���nA�p�����jVq�b�����<��iy#��P�{X��4	�۝ۧ�zI��T-orW!mPU�	o�O�@�v#�LM˰�R�jS�9w%KI#�pT���ZH|
�j�8P�E�H�㰡\�S�a-�a NB��T�Ɨc�'Ͳ���I!�Z���ޟ�������������"3����"�����?���J���{�;k���M���A��)����I�%O�`����3��nb���i����N�-^��8��7:B�Tc&s�pzz|$~F���P��B�q��w�s(F����y_��]G2��l�q�����c����p<����'���l��.rv6�W��(x=0�WT����0�8
Ά���k�� ̶���w�wT������u���������9%dcw���D��&8=��D��V�h"˄����tB��)	]!A��D|W����:�5 ��[�Sq��C�i�K�O�MZ\��|1rj}��&�Fv>aw,K���k�������G�7� 4�x֬\��Z�:��siՕ�'
w)H��=�<��miO�9p�&��&f���G��eM��W�QO�"��\�������'ڴ8C[	
�w��� ���y��Ox�#�NM^�Z*j¦��M��a��yxf�\�<v5�\X
�%j��|�0���H|��/��'alL��ҝ�E�C����� �C��N���׌�Ry�5���IP�9�H������<�>��T5��j�\P{��s��/�\.1����T�rC
*��� 1���%�ݳm]��Zq��Z&����W�`�i7�+��P
���ǥc�[`&K�;_�	��A���z����:f�Q-�����{�L���Z�{r"a��_�ۮ��n��/|�b���?I!��}�q�w7�q_N�k�~wl�8a�6�����4ލ�kB��A+�+�B`�Ǌ�V��p4��f����(�f�K��	��:rdPJ�s����J	��Q&�(]Mq�{fo��&L /^���S�J`2�<͐����:��dP|{���Ҫ���]ǆ=2��b\q�#6��k�E�7����|����&�W?)�1��w�b���X^f���o�e�KcV�Q�B���W��gO䭮��PZ���=����*�1xK{GH���������xD(�:���-ܱ�T��>�Mp�
�
�)�Y��m�H:䕈�߁ā�i��UCu�,�^ꐾ�B���<�{*����E�UG��<�`t?�g �BV��x3�;�#�����D|rA��?(O�D�Q'�{��l2��UG�s��Ӏ`����t�1A*h��ƷIڦ tۼ��y�Ǒ&ǉ�<�)jĩ��=���w��鿚���>=SP���-��V�������U�:��7m�'M}���.������e�d8�3Ǌ� ��wQnc+�E���RE6���	n���Q*S��5���O�^�����ŗ�u8��Mf��k�)����{Hgo�gt3׾�C�0�I	��\֗�j�'����,,��a�D���PKv8�@�,sDC	�_0�����!���;	'|;S^���f'e<�(��@��@�(����1W�#@gJ��-�/�4��iǅOKQX��U�X���#4N�X5f'3��~(��c@}E��
[Zz������5x��|��A�b���)*ﴙ�T�j�0����5�F�(��ޭW��@��JX ͘O�l ɳǡ-��W���_ZU>��
B!{�A2C��jȮ�jC�Q�)3t�V���y��t_p���u�-�`�onu��ŝ:��S�K�՗�c�X��{�z��Kg���C���D9���KN,�yn�ʶ�Zb7l�Sc����� ��N'd�{�H�դ3�����vf�W��<x}���|>�yYJj	
-T�{�y��b��R�	����02�k+]#S�MC���#�K(�+��ι��4�F���)F=xp�(�����J�8��e4^%u����@y��=���a�סpR�>'��v�F^ȴ��a�$�r���7�+\�����rfb3�8c�N�oL�IX'�Y��H��gX�Q��P�,5�U�Eg�K�@%���.�TSב���зG�y�r7.n!��ـ�,P�ӭ(#���|e(���V�mT���	H[��G�&�'�srW����e͐��IG'̐��<[S}��g״^����X+$+���k{E�c7�F<q�E^6�0��	yb�E��y�r�ܮ�"͕�����vD����r���*�{��~�t85u�4y��1�(_d�W`�0�Bd��c�Ѣ2� ؄�����I�ܯ�����`�9�4G�ҟ����B��5l��ZV��s��W��r>����cG�@kЯ�Rz.��녋?�9�Λ���ޞ��0�`�8�+�ꤷ����1���w�J���:k�[�'Ш]�rOo�X�`/|J����$J�o��o7��~�1� ���7H�E�/P�)�_��XJ�٬�3�Ɓ.�d�<"-���8����B�VN%�ǡUU~$x��t�͏y���T�f-��&&�	�����[���YE��<���:E0�f幏f�l}�z�������%٪��������|x䰗)�	
}���{����p0����Z	[�*7��Zi&��wᓞ�[#5��97L��e�v�P�h�a�3Ք��mHy:�IB81� Ͻ�(�w��	*\�)�טl��Y�p �d�c��g�~�,��'��;_ �k���q�,�9�Q��$��y"��2�x
����WK}��4���>����{�dN�SG�����9O=�]�CɈ���t#b=��?0�Sg�3��M=�c �KP�v�h�^�z�	�C���N�[�����։�������@���Z�I;_�-��F4p���=�-��@c  �3�P5��P �ap�݈�_$$�i��1�S��)X��u!�l�z����7���b�����(3�DUa~�E���M{Q���F���!�[�o��� |������Du�^ʦdI��{Qz�toN~R� R�]4��'�뉾��lQ.�M��UV�ԍ�Qc�@����v���M��* ���7����^G���ؾ��h�lj�܊⪵s�'���D}8@���"�G��ãe��L`j<I����|��HN��%n�ϢvE�wS���F\�}*��[= 7�A�o�h䑡a���*�B&�_tr�Ŋ8&j���W��.򥅜3��Y�I_�pj~���������+�U3u�@?l:Hz�1�d��*�P�o���Eb,���@��iqUq����4
6_��F���vp��h�1ױ�G��F;Q�h���;s�XBB �m��S��Q�)]�$�+cN4?)�P��5o+'J�W:3��k��g�	x���Ff�>��_�QOR]<I�![G�g�j������^�Ƅu( �_����Z	w���v�c�2�kpԋ%�pN���wZ�С��iZ<6���9?w���r��Nc}<�>���Ulט�Cz2f��p0IxK�^�9_�+ &cI���[n���J�`�g�(Xu�(Q0�N��E}ω��w���c��}��	��h�L��/��HB� ·.@;�W��u�h�^��5��R� t�ā�䪟��ğ�)��?�%_�-����sD�#��#���(r�8�'�hM�,?��jbĆq͍��s�$�ճ��2]���k�g�mTE��: ⌄{��=r���a�{�8�>ׁV�Ql���$�vGR2>�IzY��z��
]���@Z�d��JU�R?��ʚ�f�)�)�8�{�M�0�8%�꘬v�S� �a�ҷ3_H�Y�	���KEb�+{O�����*��^�pd�:����u<�/0�p�>���1�&7�n�vD�mS�>��QJ��L�,��a��o�ͤKꐔ����;�[E^$sH�r�o��'o֙�y{i�ó�K��H)����o�'�9��B&��r���w�H�'/!H�i�D�M��i�v���qk�l+Q����x�K3�=������k������I5N�:!)����I�@w�t�T���xY��ay�"��Vmh,h;��J�A��xdhα����T��������̙����>W�M0�U� �gawg��:W̵�8MsJ�-�
GE���1r��O��A?٠���h��W-a�7�����d����	�bY&&�Ȕ��+���}u�C7��R5��1|H+/\<2Ҹ��8 �Kq�A۴��3�P� xy_ɗU��(/}OQ3hSwO5��'M�iحv�"�R���NRb��s�7��0��)���&�x-��C��y� ��a��ܴ�&�<�DA�\u�{�������S$ ��7'���1ɱҰ�	@��w޹H�����뵀�2��,ɤ;�b����eS��e/Lm�M�P���;Ts<���@|iL���c4Ōh�k�({_u`g8�A0`�L�����y��,W�'�Jl��#P<���E�q���|���	�J�&��:�3��,Y��x,�cG��P/��/�	�pǑJ�w�E��O�A1N'俭Ŵ��|Z<�4�\��Y�@�2LM���P��t�s��nN��Y6�
�+�&�+�R�e�1���<;�	 �G��ŃP�C�\��<^�g�#����43�gl����nt*�S��n��P����5�js�f�f�aʾ�/��K�wJ�=�UD�G���d�<��
�������oN	a�fLZ�\��:N����]';����ɠ�Ll�;q_��=��u!՞�0e4�RB��R��f)�YR�|���G�Ft��le�)���f	G*�8��-�0<±����9\�{<C}�����Zѡ���&Ʈ$���~�@iqB�����0�x‴R��@����>e�=�L����X	�\̯(�ph��,B3L0Y(����1	
	��3 �B��9� �;k�A�7\�OW���`-�su!S�)�ߞ�����X�;r�!]DOqE�YN5��Ac2 v�Z�Y�Q{�Hrp�X��N8~M��&��irz��	$�\ �z�˾+n��A-on�7��t�b�邥�mtqV���d�9K��R��̘N�c����D)��e9�s����_������Q�]%��r~��1I�6�u���R�J�#���f%��߼U_��Y��{{Õ��M76	���\��b��o8*�T@!hUo�-�?�	�o�c�e��(�\꽔��Lr�۷:p��ѥ�r��ŏ��jfU����b������F������)����v�o24�R�b��(w�+oN�ے4�*���yU"Jk�[raay�E�L��c���aP%S��3C��If�u���H0C�p��Ag�$䃼w���2_-��T��Z������ �*���)x
��"{�]8� S����������f0�#ﺡA�%J���@ǞMfI��e~	���w�dR��g���^i�/d�J��	����sGgw�N����,�R��>R#�E����b�"�)��e�'ǇXv���ׂ�wB�����.��~&
��̋�=�Ǐ�<���-[�u�J�������3_^6_�b{O#�\*�\���}�
"��HSM���E������N�^�ר�a8��؛�`(�גV�%�:DD�B���S�>��nʧ@���G�x윧��Y�ʈ���XT�޹���>ݬ�Ҕd��FT��ZO�w�g"*�yj/�X��y��p7n��?)/���ilv%,���K�=�p�r%��t�a��i�_$���o�-;E��eO"gR���Q{���$��m.�O�J��X���D2�p��y�n�7�2Q:�-��
YÔ£��uT�*V?ZGp@�%0�`�˩ y�O��U�k��Q�\W{@L��ף��s��+S�}����9iKvL�	�������DYv ��I9�tD.	BlV�Gr�|l�v�˸Ѧ��=����0�ߛ�&����Qs�/�0)p�}����/o+��Lz�d��5�����HV�)�YBQ˿ōoņQ��3գz+��V�/�^�
�t�$����Vv'�Ue�U�A9y����E�?C�-ϰU<+��@F�Os~~�C|v������ZT�i9�5p�QY^�<� '�k"����jR�SE��i���/-�Fl��m'\],���^�qW;���Ш���r��%D�&W%��1�?.õN��Sϊu���������y���X�_��ð�����v�6�U��l��=�*��V�F��F���؜1��ϧ@MK�*���#�{�?t��ٸ��{�E��1;Ώ��>#N|��y��\�'I�u�_L/�U�"
�9��G{�ȅ�	�J�V�w@�i]�V°�!�-�R�t/!��j��)	��,����ͱ�k�CI�[eDvg�3x������U�lVQ�F!��]x�˜yh{$%�*�¢��V[�[0$�,X���,���H����Z�:QfWR=�1 �fu��W���[K��ic��p�k��Z�.�Ϛ;��|�´��r����r�=�Q�=Jӄ�Z��	�����>���W\J}Aŵ(<39�7�|�-t���
qW�(�Ơsk��A����d�~����B|��8�M�T�N����% �؈�Nmx:��&YIt�OD~9pΊW��q���m. ������`b\;k�L��-���s�j�����46�<�z��`�Bt:�#���@�Ҳ���ڋ��m1����Q����oT8]Ndi�7��G�?��� CFҿ����v�e)BV�qR0��N���6O�f��ZZl=3Et1�؏4���7�n�+�����ܒqWt�T��*͏��m�$r���*��Y�܏�^�|I�Ҡl�)ԝ�K5��m�-z;�}a�!�8��*F̺ND�a0���7��l��&�n��g*P�xz.�)��O�B���i��?��8�<�Y�!fέ�A2.�Sf��O]���J+�P��E4u�4E(8
����/fwJ3�9�¹hKGCA�����k��n@Q����]9�񅨽���nF����ZhR0'ܯ�y�˼��f�tDp"uβ��+��b�5q�,����N1��¾���׍&��wYv���u����h���͌�|�Y��'9�?ŏ���#P�|�N�C ��|k�a��,�*w�~k�43��񄯍�2��(t�h��t��������{%�Z�~�n��~�ㅹr-Y��~�h�������n��{h�� ��4�ܣ��g���А�%J�\��w�	$Ӳ����C��|���Kt�v��2>����6�(e������*�/`$=U���I��a��Eԅ�.�Z��cw���Y��>mx��?�c�:�Hv���p"�Q2���>���&�@��+R곖W�e�q�W�6��L�q����o����k��䎣���
���9���j@
8M7$$�� ���9��"�]�
d\�m��'e����<C\�܍��$�ݺ=-�o|����΢�*��r��NŶ��r��L�0��N07��4\�PE_�r?b^"YP06��OObE��"s��C�}���Pk��br�&�Oe:��]z�~������McBt��Q�_����gJ���m� �^����*ЩS#-?�F��$�d�0�d�LޅB��g�ҕb�;7�K����`��ĭ0�1�O;��wA=6XZ���-���#Y�Ҫ-�X��h�(��-T��p�i�Ý�n�L�b�����	HܡL:+���`�fٝ��u8����|%����7����̈́�����y^s��Xkd�I�;���c	�v��n	�t?&�
YjR�:<�`Fb���E>�{C�f �O��-#�)'��Ngy�əl�]q^�������w%�Mo;��n*Y�R9��QV��7�T:�ǬT� B�J�Py�-/%aM�}mB�[�!��g��VT/N�������-�������m)<)��� 75^:'؆jf�5ԝa�w�0j`]��Sg�jV�G�m�Y�������^s˗=i�����β޹�/S'�x�-,&���!�_�+s[�fq]�{Ő�Ӯ1�Ez��b2?����+����	A�L�m^1�3@�)2�v��w)m�b�%]ݖ=�y��*������1w���W�x%d�w�zƭ�'q�HMW!!�"�So-� ˸�}��o8qf�Ȣ�fi���:�N8���s��A(?b8�Yv���SD*f�e��hu[<���C�6�-7�i1�>�We �6��8t �Z ��Ӄ*0���Y�K59D_����+�p����
tJ�<�/QK���ʓ���n
+m�$3o�Ϸ�����(;u~��@e����
A����TG2�"x�b��l�B5�y�ǓI�/�o|�����'�XD�s��,8�v��}Čfo_T�+��V�P���������o�b �GC�y���,�m%��G/���ʆ+�6�͆�;s�fb[�/*�5���ܢ�>ʔ	j�N����e��,VzO{�ڳA>\i�3Nf����G���5�~k�����kY1ʎI�O�\93,�N�X�VA,q ::�4��f
){�h�DM�MWA�?y�q�"|�e�*3�"%�_u:~)Pf�{Uz�|sT�Ux{Z��T��0��{GCȬ|B� �`�gyq���	���b�O2l��CwF"�����ꇾ���ZE�=h>�6x�'���vs���� vȊs4������H�ɼl���x-���!۲I�wœ�t��wJm�|>&���~B����0X������=כ�V4��<D�HEE�<�j���)R8��������,�ñ�ڬ�jCf�� ����M�0�t䳟��ĹO:&!����x���դD�F���IN��tp�� 1;���ه�,Ҽ-�%�Uf� Y�}���BWC�,��u����X�JW�[i��+1n�ѫ:�$	 Z�ZᴞI�B庵�Y�Ga�LW�؞�L<3˝�vG>�[��D��J���T{G�����=~��I`#��ʫ�����,[�����7�?� iX�g*��EX�������������ԴT��bm<愓�=�Kk����`������~.��;�(>i�&�yZ�x�+]�#�ɧxMbguWg RN��M�7��M��pVt�A�XeO�5���^1�%~CϞ.���֯��L�������1����3�p����@c�a(_�5�z>=���;�6�`>Deop<�&{��v��OT��ڬ��u~��D���9��ۘܲ��3�G�V!�K�	<R�^p�)�|����R+N�6�|��P� <">s�v��F�yb����k`J6�͡;������S�����T����7Y����d���D�WeA �ͳ�щ���Z%�i��3���3=�6ڵ�K7W,�00c
��>s��A)��"Xn w�ׁ?Aʕp���yt���?�7���Fd�wE���؆iay��Ċ��m�\�Pi`�}���3�t�4
�7E-�Ģ�c������$0��4������aǓ����"�@捃�ou�@x���/m�$J���,e������#/pt��.���uO�#�j���h�b��<����s�	�9m����2�" �"��R"�l%���Q�
�٥��?�$"5S�X�����u�/IZNb��%�i�ӧ�����{��ǝq��"a�����qj5u�gBoѵ+ixУ������1������s�8�oL�K�����+�����ʯ���1������ْ'���݂��|ye��
 |��!��_�L�g����g�<�zG�df_SD�^AS@U|	Z�'yٷ�t�|p#
7���pM��̳�& �c���nJ������M	 �S��m���ڈ��sF��-M�<��{�`�Ȉ�~��qK���e���� 	EA/���gɬ;z	a��^a��]�/��ƕ1o��&~���}��%�ߪ@��61Q0=QՑ�����5O/Y��
�Q!b���Qu$L�L�$/�݂�W���5h̺Xص0��nC��tz�R�RgA�v����D{/�5	DK�fYǔ�=����L�2��W��?ܥr{2��Y�R�is�-H��g�Q�}f9�8µt��Iw�4����H6ؒnk�U�F��N�}2}�*�C�s�ƕngk��D q̼�A����0'��3��X�(�`�4s��˲x..]�j�>`۵�܏l��ZvKk�*d�!"O�'Ν��0�Ӊ{�ܦm芴�Fz_�. o��o�����.+�:�D�zjAK8;�.�tl���Hm̞VP}"�tz�=N�����^����%$���{R�1�ؚw�Ȏ	io�����s?�y�[{;�q����M� Xp*��VBs=M�wA[���ܰ�=�`	��1�(�%�_�d����%?���b?g�_8 )�5�{�mٷ��xu�4V���SN޷'�im�?(���O���mۃ�&@�ݒNL����D%��Ϧ9i���!A�����	�W�N��X;���t����+@(�������E��:�03�'h�e�8����8����c~A�GA�@ˆ3��
u�n�&&3И�4��cCJ���V= r�}`�@I#�P�#�%����v��p����
��Aߞ���� S)A_�O� ��(~<� ���B�ȿ0"
)j�
��3a�����e\��#m
�+6�(d,�l!*{aɎ�4�'����{v&Zx&���n�y.֬zӹ�{̈́6-w �ґ���z�������F, �'(*[�`���"I+�a�-9�5q��^*�o�{�r�p�֭����腢M�TM	�r��crf����������6<��D��{�6u�V&ޤڼ�<Uª-��� �;�������A�*�W��]t���g��b��-�)