��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#�?�l��Z�F3~�Qp|��:��pIۄ�d�
��&��Ađĺ�M�����2�m��ahdH��I�*2L6cB��H��&�a&�sۘJ%�b��T�f�%�Kz�-�����DU���<B �����r3�)m���g|��jC(��:���t`��d���\)�b��Su��ʹ��ƵV�%�KhɆ�#�*�u�����Y�wI���h��"�h	xɑ���_�KOp	m�!C�(؋�	!{V�GOf���W*q]�؟�r��b���PM$�g�S�%��6�7�`]]�974���X���Hi�����N���7m����YS�v\}����B�AfvΓx�o.�$�dU��% �FF��}�-�Q|�k�cc�I���5�N(<s��%�L����Í2�n�|���"˦A��z2��m^�c�:G�iEJO>�i[�� �hm:nG�t`����e�8�L��.�f(����;���GV_�����A�$����d9���P�s��'��B>Y��<[R?����R׃'��L �I��uAb������L*L����/X����
�C���Й���iX/*�����������W��T�Ymg�k<$9D���&y�S���x��/m���H�\wR�#�Z�3��&�KԖ�̰�fzL(��~J)��
qV+�)є�c5+����#ڌ�d�i+�+����<&�Q=�&S��O�7��T�D�z�)���u[m.���F�>L����\�c;�
������|!�J2RZ���>�r��_��f����;M��x�F; p�3�pC�ƍ�p�ȸ>)ysLL��s3�(~����'������LONh(������;���v���s�P�Q��9���%lx.�eaUj���� ӛ��!|s�\9m�?���o�����G�m���ϣ�<�����[�6ߪS��\w�������V�rV������ oRq8�!�0�~Ӛ!�M����*m�W��o�&\݂f��5G�!�z|�q�Pb�`|֌�A >�2js�Qǈ�!�-Xq�ݾ6�ˆk���DY/in��S6!9/q�dl�q��6Vd�tތ N�����j�3T�qzA:"�B���#J�k�;4a�����ϨV��$��j�<������]YF6�`��Ī9E�V��V���NcuۆY�)=5t�N�j����&��-����a�`�;E-�)ORЧ���/��-�T�h�6�P�Lߓ�(o�rw&T�hUZ]:���bv�pTV��&I'��/�^\B�,���y�wm�I����_�P�
�l�n3�5�0p�O�Fm��l
m��^U�g�2�K��Ƶ����CV��ř�J�q�[Bk.Y���-%8�[}��*�]�aX\#\���k<ʯ���"��]_OKSh p���nz(<n�)N��ƿ��!a�������I���ܛ
�#�5�D�hv)����
�j���Y�����`��
S��Q��l���<��e�%���3���(���)Ԩb��cHO���iC������t_��q�ۄD'�kVA>�;��\П���I>�C������������r��o:uQ�8��!�Ԏ�������A�����|�ț�A��$��m������ɮ�k�-����A�V���bE{Ueݖ��5ȵ�ח/��?Uq �����26��Q6�/��>���P%rB��JS�1���X��4�ۏ�e�P�W���Û���*R��d%�y��SP9X����^o$���[0�l�PW	 K�x��k���\�E�f�7�lcj�v0a�JW$��(
�;�\����ֹ�/=�@��!���j-����(� i;o���uG����l��y8=���@Yd�s��8/����8��@Ӭ"6|�uJm�kɵ��p°��ƽq�{�7�b�P�L�Xh"�Q6�{�鿆�=f����'�58��4�st�8d�_E�4uO;d�"���t)�#�w-r�M���N�}� (� J������afa�T�Dc�s�(X<or龏�Y�9v�|����p��.�;��b|�L�9��~[�/_݂���s�#���cf-��&7��"A�¿ ��,bF�EGw�G8�Ķl ���w��p�i�p������������k�
����� p;�k�~u�9eJA���ߩ0o��.P��f��a�rј��פE�G &�'�&���T�F1]S��iS!�c���@@v�AZ��`yNP�y�[���?���7��@T��mI�-	KP/�U�tƧ����ԍ�͞v��|����x�b=�A����g4�kB�\��b;�0Ĳ�z,�zα^�����z.�wg��=�/�6��AW�c/���	~�e�_P5%&&��p>�4�̖WlwX�Z�E��"|���;&���g�ZA�XB����h�����8 ��O�0���;�6[*��Q���u��v�萄KI��du�����R����DXxC4[N*�7���k��{�Ir�	c+�tu+������.����o��1��&�~<26����S��5�rP�d�^��'��ë1��@c�;�ػ:�|�� 	�9?��Ҿ��W�Ӿ���F�a���Բ��K��<���u�!��=��+5��P��'�b�,%T�ةi�}燘Y#�?������0�҉v�w<���V85���6�Fκ5Ė��r]gR.j���%��ߺ���kN�e��+��O���܌C�"� z�N�*6�Ie?"�,�l�J��'J-$o|E$�����<V�ۜԑn^��_!�__u�w��e��a����&E��]�:G��Y�jh��&�"2��<�c��0RG�T;�������A��?1c��\��w��d\�,D�����
��l�2�q[��Q��Ibd~*�:���j)1�e ��]��\�~gK��"�����z�N� �76�t����o��笩�4s�β��qV�:��Ԅ��R*��}�\󘶣��3����9���Z�	��k��o���Rȧ�xwY�b�3��t>R�C������ol���BrQ`�����An=������տ��,�k�3��vu��EX���v2�޽Rΐ?�Z�k�Kgs]4L��������>��m�q�]{�t��y�m�5�8aڴ���֣����`�I��`��̘y-Z��r�V���[�/��hAw���z:Cu��a�U�Z����p������Zn��e�fw��;(ĴY%��!"�.���M�a%��\	 odɔ��^��y)��G�� �m_��B�,�F'(��Wi?q�q�/�ou1��"�y�v�SX�~y.E'��oY*ֲ��r����X���Wc`63��������!~�1
�hc`,T{��Y�zA�n'Sb&Q�Nr��ʗ��N�R>�ڵ!�:���|� �2�۵]AϤ#a�ڠ�S_�ޔ�SLGscѶ�'�(s"v��ߥ9��+��G.����0��J�Dڱi��r�i'� e�^<F���S׏��B9��B!R��n�ћO.x7vx�>��.)���@Oy5���G��V�� � ��6��DR���������wkɘ�}:���~�.�P$��V���/$��I����'H�b��#�y�� #5"(tI����#������6�ǥ-�RG2POsV?�ߒ��<������\`⌛��Q�@�~h};�H ����%E��ix��"�ш&�`��o���� w)P��o�/��:��ЌW!WԤ�� J#ox���%��6��+�߳�ӭx���

4Pwߢ�5����*f̃<�Pj���+:��8��1J/��?79��I�œ���E�V�8�R\�Se�t�cT\X�I�Z��f��|i�B�\�Q����v��T?0F�O���3�A���)ћ-}M���!��ǡ*oȝ>�ge'����<��9�kI?���Kw#ʠ;1|�r5,�XVeLt�n��v�i�Ċ�1����{����h7�l��u}�$��چ�#�阋>8-�ށ��|��M���4ҡe��w��;=���V�锏�l�[���U��ABª�_�*��	e�G[Ӆ�#\��i�R�%��K�Ƃ&s�~��)1���n��AI��s�%?��4�}�������*@@�I/����?��Z=�!Sn�������L�'�u��k\F7�y�I��~��`�5B���F�
1?ӸbՖ�?!^f��t0��%��R?h�P�S�^���*��
#?-�m�������#���d@��ؘU��f�&��w{�<���q�֬$�2N����A0�%�a�F���]e�X��c��������'
��z��BWv2H�,f�&��@%5���ڼ|����?�GK�;�\���&f�n琚���d�dB;H<�,e��P%�<�[�=2�����έ�+��_>ߗ8�*� ��xP��Ɗjx���?���ɼkRF������tᎈ�:H��5��Λf�EI�A�ƣ߫yk���yT\�.j���k���tY��g��vy����ղ1+���2�)��d�C����Ǹ�X�h]�#S�o���ҡ�
� ��cǞj=���ܼ�t�=Џ�#WZ�3u[�lF 
�X�)ŧ����.�����
Ro�����Q�3<5
9V�r��)�6�1��y��臎�[|U���u��Z�Σ�"���>ת�dd?�?�)�3J�<A�����/ݞs+�k�ϕX��_�RI|�q�:d?� 5tg���++�/�``�X�(���
��8:8hC��'�v�Gc�H��,��sc�� -s���63a��kf�[f�f��� ,y�4�V��gn��Ւ�!�@'ڎ;��7 �2���<�Eb'�H����	S��)6�p�xvʓ�ǲ|��{5��OoA��� �=��PqQ�hF-���e��M��b @������r��o'�ȇ��X��vÆ{,�<�0$D��{�Y��B��+�Qv���v�c�>�č��ru֮N���߱�Ww>(��)�d	
p|v��m�C�
�܅�t�f{�]��&�P�H�3~AS!���k�7�s	��J%�3�H/QX�S/�m,9@�.�0yc�/����:�+h������<�!��5����̌9��W��}��큩
!r4�Uպ��ٜ� c6y�ڿ��+Z���0V�x"'�@�"c�W��cI�}���f�t ��`����C�� ]y�j`�/ԫ�V��&��tzn�n���nO�G	���Xw�\��*\���x�H�S�������z��<�kV�u�K��ٮ�����*����#��6��:���r�ȓ�(�������ޯl���-�Ѽ��dȻ�A�
v��F��2�G㖯�G�}XAc�3�)X~������*�������f����}d�,����Vp���o-�FW��l~������5����ʁ�Y35�lj����bT������ ��ʤ��P�Yv�8A���|���Lt��w���hҐ|�Bs��X���V���!���:�j�k��,_6�ى#���0�(�� �v��[�z�,�H"��>��PX��8Ug��Q�>Մv�Sč%��}ͧg�(�D���(�j�|�F��b�u!��l�xܱ�-Z�O�t����x���r���sZ��XS�+��V2@�ú�C������n:�jޙ��3�י���6�b>f����F��=l)����q��ą��R1�l� �s7*�Sn��Um�,���k�U� ��H.z�,�ᙒ��cI]vuI�cu���̇��"�I�=�BQjA{m��KR���?�џ�+dT��	h�@5��[2q缭��J�8}��YX�F�)R�['`�U�6M��%P(�o]�
��C�J��͔a�.���4��f�_�6j�ʻ@7i�8�`n�lf�E���t�ϒ<�[{�V�Ў���Ac:ՐCc�u1[��F�9r���N�.���=�{�$ϴ&����Ә��� k$���h�	�~�	V+�2���5c�B���sq-��(	�4�T�Uf4p�c}�l/Rr���W��3(�$��sI�g�"t��c~s�� ������F0kR�|�w�?���e�����W7a��n�A%4m���ߚL3��!�+�͢�;�r]��/��5.��)�ab���ѓ��&��{؎�,�ޜ/���Y���_
k�=�*a�1��?�p���G��4:�q�(L`I�Nl�L�<�&鰶 ���8~����9�T=L���1��
f�L���Ш?�3Y���9�;�'k�\����y�������R3LZ�z̕W�2ߟ\+5��o��`���j��R(7�wV���޺��!���G����}j%,�CP:͗gy
�0�3!q9Ǳ6Ƅ"+��8P|큳�12�el�oV0#���ć ��Qԯ��7?NK����謹�zDe��f3g�SiKyU��wC��r�C�/��dD�&�Boݡ�X�U�L�=����Cf��H�qp�C��N,&u�!f���gdI��_�e��it��ػ��x@T�54�Jj��+7L�C��$J��s��s\]�+kN���1�،�2��&�g�׸�׹&�^��RҍlR%�]rW�a!) ͝}��Ͷc����-��m7;"zh�[����Ry�8a��NKƩ��BƜ����g������e�(Z�%O/�"��E�~�~np���u�m�A�w��8����mG�:I·U������p��r�@[�u�%�W�!�d�U9���f���"�kk�Pi.); ������b�s�^�F�<�����-
�wֲ��ٷ�&���C���xn�Z�Q�̼o���ʏ�T�Yۜo�h���z�B7�$���Ԁ ,<���a �A��&3�$
�GL�ԕ�Xj�=�ہ1�/���woV�<�]���h��q�4lG�����!WC9�@^�
/Jj��`2@�6�6�X1��V��ũ�k�Uw*
�����簧�����e���}T���l�@��L���e��׏Y�b����ea�dpU�1�9W]>�D��/n�	EC䅟��p+�����<<���C�bʹ�V踼2D��I�	o�/�Y1��dkt���g�3�j�2Q�������y�l��Z$�OD�6����	dL��(Y�%�2G����ќ�	� d߱i�_�E@r	?�>�G%�U��A�Ӷ.bUd�
p'T7��gQ+��E�$-��?���Gl���X�E�8���}?�DXJ�`F�&)��a�� �����e�����\��p9���S�nI׏lm���0�ϰ���FKJ��'�8�f�M���rM(�4�I,�-�XLW`'o�)�!�У48645Ӂ�8��-Ii5��	8�e��i�+R�i^S�ۀ ��iz�@*R���A8�u�L� ����|�����ً���s�|d�̌��MTs��p�RЬ4�H���v��.W���i�<@Uc(�������"
�x9����ɷZ�Z#'6gs"�]�P�D��S�k���m��e��W[,3�n�jOn��U9���P���/�b�<2*�iy����92"�d������w�LH�-NMs���v�7�Fh헥ݲ�z©�Aϧ�ޒ�su{؄���\�z�&F�2It�<k����-�<�0�>�}Q���fz�`�x?p)�[�!xi�;�H�nu ؋���}��?خVn�j���q�y�փ�a.|2������̫:""9�ff�"���Oj��0��9�?'YB�F�s<:O==İ���ԝh�J���<��l��[V4w�~�:K�g�Ƅ�?9�2��0�q�%����Nd%�QI��D+4o"�<B��'�&8{j�eU:%.��e���x):Q�F(�hޅ�v �<>d��P����y�o֫��5��$��.�o4�ߜP� %"#7b~��h�ۺ�C��RM���N\C���h3i�*����/e���"����:�*Xx���W��(�G6�aLqM����)��H�I+�lEdW�i����=�_��� ����_���$D������4��wJ�(�vS=�	�t�L&@yP�������/c��ۯ����QD�8�z�dsl:Y�{���lM�6�á�c�ؕ'>h��eN��Z� �uG�n2�s=��`��i�(��c���2��BH'oF�=\0@�s������cz��D�k9Hhg�1�%�ꢤUp꺼�X�w LK���]ZY	HDV_COt��7�����*��[8�v�c�e�vG�<vi�!��ߺ����@�c��N�����$U�0�F�����q�t��S���9Եµ#Y�c�En�9��eqrX=�E�[&2��<�O�+i�o��>���U���?�<n��'�y_	�F�4��t��L#l1^�xO3Z7����1����q����{�'ko�f�L�v�k
� ��
�)(��w�֒B�f�O_�&i;:�tj��1�[�4�曲���"�u7�M��h&��q �����L�2��o9�X`d��>�H��O2�s�E��?�4z�+�M��h���q���/ ���P�:��#���h4V*�'�@�u��&� �m҄�����	R��w�E�*&6��s�9n��_��t����&d���Nf:��br���z�t�%�C�8�&I*Ps�Z;�W��3������G2
C�*J|�R�':5�(�M)_=����X6;Bv�sc#i_~�/���)�s}匤�!�P���3z+�O ��'�l��gI�e1�q�@�<P�v�	�XJa#$��0�ѨI��.|�n���@�e>�p�k,;_:B^�-�P��i��ԭ��O�{`