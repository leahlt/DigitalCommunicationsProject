��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P����z��{}H���_Q�hФ���]xy�0�|s��9߼L���حe=�3�����Uh=8G%�t���n�4��D�cm��zۜq�a��?w}HC�#u¨�`�L�Cަg
WS�1f�k��Z�WЁ��ehg�+ݖ��F�	Y���җ��2)W��Á$��%��-�B���C|;\�z�8����P�����`��:���\���c��E�14�QC4��l���&�d�2]JQOmF3�����A�-��fIF�_a�,s2`5�A��	A+�2�F�}�Q���y�4�k`
��p��]��y$gk;�#��)Y�$D>�I��d��2��'c��v-�� I����)1֑�_F�'���B!��v�J����e��e=#p���G��(_�Qh���,>FaM[�c�u�tm u�8�R�����o��&I%b|��g�C��k8<�<��h����+��1�n��x���eAe�kXn;Θ|2N`L��9��F
���gV���~!p���f�p��m�t����ǌ��b�l����aZ��k-��{CPK�g��Q��FM�+$��fp����қ�)����Ɖ�X�ё)�L�ֵ��Pxȧ0��55Xs�a�ýݯt�#���?������@%��d��L���Kù�)��2%�^�C�'o��ݷc�C��Ol�W>j��Ӣ#S�)-/��\�l�mV����Y����w�_F�:��]��a���!�_��r�o���w.J���z�����:W�<�^����AxЯ�X�%����wk�A���?�԰V�5�?�|TS��>�}�aL�,v #1
+����6w��Ѭ5r)f�z�Q��&^O���e	�#E-F��Z��3�L0�<��x��=�1�t�����sv1H��"����G?�֨":|x�_�sMH%w_+n�����c�2>?f�F���W�G�!9��9+ڧ���'��h��uڇ�!�ΰ����l.�Oϻ�U�"��V���[�7pbw�f�Z�.[�H�.�[A-�Q��&U��)c;*���S�}�.)����m+�z�V�&�ˁ��ۿ봴�d�#���}t�e�嘥��d�E����Gu�}��	G��HH��ml��0�V����fH�> ۉ���+B�D.�h��H%..�p�U��E4ֶv�Q�1��|���8�`�R���:�}V�y]2j$�g�\m�U[��d!�c�(�C�T�8�*�X�/�o�OڈQ�ݚ��`���H0?�!}u�|�`2�~DS�^ȡ�]*�N�����rMu�m$�`��S�N��Ar"�_������ L�,�N�Es�,Ck_5�h�O����Io��*_�"s�*Sq�L��^����Y��)K7	��#�	�L�m�M#\�2L٘cn�XF��������-��;�!���k;�\z�O%d"�/�~���gU��"�{\;����d�?�c��|�m���w$�_Q��e>5�c�z�ݒ?� �'�6uB�f)̱�'�p����	�������-栗���,���/ߌ�'u9�"B�E��\>x�E��"�u����6X�`���r"_���0��x�:~֓��Eɲ�[Y1����{.+*�>����"�DF�{y~'{���g��r߾���R����}�� ����ޑ�D�τ�Tas3���ԏ�wkAw�?�D���R����Lw�����'Kg�CZ�"�T�Ŕ��/��0����7��Z큚 ]��~����ۺ�3��AH���3l��'#�+�C��A�t���������#�����k�.�=�V���Mo�����w���g��Bsd9�~��-��0Wd��YO_�K@S�"E''�jfA����0�h*t���)ye��Sc��%�C�7�(��`��6<lgj�����A��ѣ����(��#����jg��|5�ZY�&���b�"{���14hÅqЈM�@����8��L��
���0'J.iѕ����5�B
���.�$�ĊI!<����5�����x	0fRZ.�W���	ƚ!���ۖR�{�k�(0�� S�w�����
���Ө�ӧ%�dY���S�=F�D �e�oث�8,֝�j1� v�+:� ed���u����J�d���]�p�%y��[������JD9��T�٤@�{%�)�&��vk��~�iy�e7C ¥j�sek�=i�bZ'��Qݘ7eILDn򊹝3��j`I�ڂt�K��=��4o�`D����²?����<�4�pR�ClF�E�H�<�E�ԯ�x���{;�}�ܷT�K�?��xXT�oh��.�Ɉ�+Q�֦�"�!<o�`�:�v2��2���ꯋ�E'�,-�.H��R��L6���|��g|���ͳ����`�a�֛-�0n�R�oC�,�*�^������� ��0v{I� M��m��0�Ni�E�
��+��Y��X��tP�p��$��+��M��\�v3|��ύ����_�����n�hI�T��}�5��H!L���!H�[N�l��_�2P�'��!m�WӊI��:��M[8�u�U($1qF\��39;X�n(DE��Ic֭��턖x�FS&5�0��%n�9��{R�?���-shs.��X����5��0+â�3���FL2�O�v�ӏ?&�~]M����c]��B�F�B7�5��I�o��T���Sd�f�n�1{��PXL�����S�E�%����Ȧo��`3�p8��<��]�w��a�