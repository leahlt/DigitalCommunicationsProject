��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P����z��{}H���_Q�hФ���]xy�0�|s��9߼L���حe=�3�����Uh=8G%�t���n�4��D�cm��zۜq�a��?w}HC�#u¨�`�L�Cަg
WS�1f�k��Z�WЁ��ehg�+ݖ��F�	Y���җ��2)W��Á$��%��-�B���C|;\�z�8����P�����`��:���\���c��E�14�QC4��l���&�d�2]JQOmF^����^�Se��j=o���]��+I;��l$P\6��X�u6��fK5��\��<�Ŭd�sz��bVWya�b�+ ���j�͜��#@��.�+�9n8#�*������0@��\�'�x8�qȉ���f�O=�*���C�)kB�D����{��l����?l���8���bj���qU�DsV���dKϝ�ro��i�4��3�Ͳ�DGlS�W#�F��� u��� p\@G��.�/ʰw�[�
/&���Nԣ��|B/�3t��Xb���Ȏ���H�Z��;��ގ�1�\�yʞ�/��설v>����+�I��`˕jV���|^i����1	7`�?5Lo�Q�;1��2�sҮ��z�
$È�-'�O��iX�������~0Ru��r�U�DnZ���sR,�5^��T��&�U�����`;6p���v`�6t;'���䅄�*�. ~f�d��c�5� �$�7k������w\;��4Ɔn1A��y��QĸU���'l���K��@{!b��E�a�3��sH�kڀ½CN�ŉ�Q�̷�k�M�!�$j�Wȑ���,��i��:��@�ele�	p|�4^G�<φ.�O��.�:dE�Òظ��n6bW��j���X�� �`+��>f�	_H�{�	��0�?�jtߑR�D���P������L�w�{�$p���]¾52�Գr�+���P{�#B�}MZ).H���:̉�sË䁉^��� ,X��P)ז~���(�EJ�(�T��Ŋ^d��Aa
�:Ȇ�&�qBh
�wb-�;l��?l�����f�6K"�r�����=!)դ�=���G?ƚ��K���}�Z1�B����"X�S�%à_����_�P���l��j�����Gw�]y�&�\U#��h��� )��;:�k;?#���肞H���/�}�k���F΂4Ś��P�t��g>@D"�^Ad�+�CgV�ogD��qx����U���ͯ��N�'�1��LY}�w�>��o�=�{䎝����Rl=�="��v<8w�3�3[��+��=�/�H��a����0� U�O�M�c#O��+߰UD�`�@��*�W�D�`�>�P]�l؋:X�V~�UY|�C��]��E� ���}d���[��e�K�n��,'�9&�Q���yl4�b*������V��WG���A�������L�=�qK�D<3��O��|_A� ��� aut	N��L4�i�W(�a?������`�]@�\�g�ye��x�ܖ�A��7# K���H�}��,�E�:Id?��^ňt�P���Zx.!�K��|��W�}]��]C�j����ܱv0{h�n�+��� ���O���k�,Iy*A�f���!\��� j/��c!�##������]7����S.����C;�Q�]�Q�#eor��2�~��/q��~�z���!Ԧ~�˼���b�q�_
DFd���r �ʫH4��2U� ��/Nr�F�[�G�=���,BXaAq�a�;i����1$��kZq���s�Vi/sHd	M�m.��t!0&D�bޖ���}�C�ܷ�Far~�w|�fG}{�eeMk�l�?�O��n�V��<��4v� �2	�5ъh+��cD��iX��z-���F��5L��c�r�P�F�Zʱ��=�\M�'r ��#��䤜�GbZLn��bh:�J�63.k���-�4�����F�WTe��,�e@��Z�A���o��N�e@i`�����9o��|���BN�;�,�9����N�2�:�+��+p���@ʿ�W��6h����׉ϻ�-Lҩ��&ˠ���I�^eqJ���Q�+3+L�5��˙�4�Uͯ���Rr������;� \0�W�ԩ�����YŚ��l���8�H�n[�df��QuzD���-��%��dy��/�Đ�s�A��*�e��osf�c�nZ�D<$=��V]�nbm��I�ҧ�x�D�������7�5�b���y�1���$�{.e`_2"j�@��M?=ޭ��6"�*oN{��-~sĐ�X�r`] ���f�ti��Z > Tc�@��I>�N�\A�DS��ӗ;J�p)yb��x/��3"t�Fd�e����+��l�CC�"����;���.��?�X�|�"����Z�ʑ~���ݕ�S��M��i�3�HZD�hU?$���J�n��w�@��\G��j�����em��������Vk��������OqZ[Xl��=��|b��o��dI=8�Y�0�I����r<�P֙1·�Q�+j�6	�:.'�k /^�t���D��D�|�@U��ʹ�&Vȯ�Gz�&������&#+f�l�?��oPny�!a0�D ��|ݧ�<�Ђ�M����v�㙝D�F/�b&�4/����q�9��BE.ZEUԋ�ǭ���<���3�;�:�I��d��Fڤ�8�=�:ԩ��fԱ�æ���� ��S�GN69+�ƚ��u��^.a_5?�-n�ȥs�;�(�CI�J�,�/����z(Π�