library ieee;
use ieee.std_logic_1164.all;

package bch_enc_package is

constant CODE_LENGTH_N    : natural := 8784;
constant MESSAGE_LENGTH_K : natural := 8224;
constant PARITY_LENGTH    : natural := 560;
constant DATA_WIDTH       : natural := 8;

constant POLY_COEF : std_logic_vector(PARITY_LENGTH downto 0) := "111000000011111111000100110110001101000001101110001011101100101100110000110011111001100101101000001001001011001110101010011110110110111101001110101001111100100111111010100100111111011110001010011101111101100001111110101010011100110010001010110101000001011001100110110010010010101010010100010000000001100000100011101111101111011100011111100110011100010100101100111101100010111111010001000010000101011111110001011101111110111111010111011010010010001001101111100110001010011011010010100000111011000101011011100100100101000000000001010011100111011110010110111000001";
type lfsr_coef_type is array (0 to DATA_WIDTH, PARITY_LENGTH downto 1) of std_logic;
type lfsr_input_coef_type is array (0 to DATA_WIDTH, DATA_WIDTH - 1 downto 0) of std_logic;

constant LFSR_COEF : lfsr_coef_type := (
                                        "10000011101101001111011100111001010000000000010100100100111011010100011011100000101001011011001010001100111110110010001001001011011101011111101111110111010001111111010100001000010001011111101000110111100110100101000111001100111111000111011110111110111000100000110000000001000101001010101001001001101100110011010000010101101010001001100111001010101111110000110111110111001010001111011111100100101011111100100111110010101110010111101101101111001010101110011010010010000010110100110011111001100001100110100110111010001110110000010110001101100100011111111000000011",
                                        "11000010011011101000110010100101111000000000011110110110100110111110010110010000111101110110101111001010100001101011001101101110110011110000011000001100111001000000111110001100011001110000011100101100010101110111100100101010100000100100110001100001100100110000101000000001100111101111111101101101011010101010111000011111011111001101010100101111111000001000101100001100101111001000110000010110111110000010110100001011111001011100011011011000101111111001010111011011000011101110101010000101010001010101110101100111001001101000011101001011010110010000000100000010",
                                        "01100001001101110100011001010010111100000000001111011011010011011111001011001000011110111011010111100101010000110101100110110111011001111000001100000110011100100000011111000110001100111000001110010110001010111011110010010101010000010010011000110000110010011000010100000000110011110111111110110110101101010101011100001111101111100110101010010111111100000100010110000110010111100100011000001011011111000001011010000101111100101110001101101100010111111100101011101101100001110111010101000010101000101010111010110011100100110100001110100101101011001000000010000001",
                                        "10110011001011110101010000010000001110000000010011001001010010111011111110000100100110000110100001111110010110101000111010010000110001100011101001110100011111101111011011101011010111000011101111111100100011111000111110000110010111001110010010100110100001101100111010000001011100110001010110010010111010011001111110010010011101111010110010000001010001110010111100110100000001111101010011100001000100011100001010110000010000000000101011011001000001010000001111100100110010001111011001011000110101110011111011100011111100101010010001011111010001111011111001000011",
                                        "11011010001000110101110100110001010111000000011101000000010010001001100100100010111010011000011010110011110101100110010100000011000101101110011011001101011110001000111001111101111010111110011111001001110111011001011000001111110100100000010111101101101000010110101101000001101011010010000010000000110001111111101111011100100100110100111110001010000111001001101001101101001010110001110110010100001001110010100010101010100110010111111000000011101010000110011101100000011011110011011111010101111011011111011011001011110000100101011110100010001100100010000100100010",
                                        "01101101000100011010111010011000101011100000001110100000001001000100110010010001011101001100001101011001111010110011001010000001100010110111001101100110101111000100011100111110111101011111001111100100111011101100101100000111111010010000001011110110110100001011010110100000110101101001000001000000011000111111110111101110010010011010011111000101000011100100110100110110100101011000111011001010000100111001010001010101010011001011111100000001110101000011001110110000001101111001101111101010111101101111101101100101111000010010101111010001000110010001000010010001",
                                        "10110101001111000010000001110101000101110000010011110100111111110110000010101000000111111101001100100000000011101011101100001011101100000100001001000100000110011101011010010111001111110000001111000101111011010011010001001111000010001111011011000101100010100101011011010001011111111110001001101001100000101100101011100010100011000100101000101000001110000010101101101100011000100011000010000001101001100000001111011000000111110010010011101111110000001111111101001010000100001000000100001100111111010001010000001000110010111001000001100101000111010111011001001011",
                                        "11011001001010101110011100000011110010111000011101011110100100101111011010110100101010100101101100011100111111000111111111001110101011011101101011010101010010110001111001000011110110100111101111010101011011001100101111101011011110000000110011011100001001110010011101101001101010110101101101111101011100100101000101100100111011101011110011011110101000110001100001000001000110011110111110100100011111001100100000011110101101101110100100011000110010101001100100110111000000110000110001111111111110001110001110111110010111101100110110111111000111110100010100100110",
                                        "11011001001010101110011100000011110010111000011101011110100100101111011010110100101010100101101100011100111111000111111111001110101011011101101011010101010010110001111001000011110110100111101111010101011011001100101111101011011110000000110011011100001001110010011101101001101010110101101101111101011100100101000101100100111011101011110011011110101000110001100001000001000110011110111110100100011111001100100000011110101101101110100100011000110010101001100100110111000000110000110001111111111110001110001110111110010111101100110110111111000111110100010100100110");

constant LFSR_INPUT_COEF : lfsr_input_coef_type := (
                                        "00000000",
                                        "00000001",
                                        "00000010",
                                        "00000101",
                                        "00001011",
                                        "00010110",
                                        "00101101",
                                        "01011011",
                                        "01011011");

constant LFSR_OUTPUT_COEF : lfsr_input_coef_type := (
                                        "00000000",
                                        "00000001",
                                        "00000011",
                                        "00000110",
                                        "00001100",
                                        "00011000",
                                        "00110000",
                                        "01100000",
                                        "01100000");

FUNCTION log2_function (constant in_data : positive) return natural;

end bch_enc_package;

package body bch_enc_package is

  -- log2 function
  FUNCTION log2_function
  (constant in_data : positive)
  return natural IS
    variable temp    : integer := in_data;
    variable ret_val : integer := 0;
  begin 

    while temp > 1 loop
      ret_val := ret_val + 1;
      temp    := temp / 2;
    end loop;

    return ret_val;
  END log2_function;

end bch_enc_package;
