��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P�Su5V��RFpg�a� (����a�	���D`�~�CLD�|��<�
�.K{���;�Mc��2ͲX��
��g�T�1�mc�-��f�8+;"�۔���[2�1� �i$ɥo>	@T/?Ur��%�I r��������zCpm���`r�3v}�sk�U�Ԯ|�n?v�M�F�=Y]P�N��6l$3����0��yX�T�����6��y�(Ĥ%���,�vW}��	��U�%ǲ@��5ȐZ[�Y:�|w�~�l{IљRoi����(K�H$A���y�"�UNқ,]�6�"��&c��|ťo��݇�A���ϛ��b���;��K h7Cɸ(��A��Wl��0m[�uBN0�8� ۫O{�� �Y���RJL�Z�if�����\"����$l��vM�w��hL��1K�3��T,{�u�����^sl�2��1�!JԤB��}[@�Z*π���=}X��$n�ޣۥuKUVB���_4$�R�'԰��F�oH������4��y� ��Q�>�*�}8��}2]7_��=v;�rQ���_l��Yp��Ȧ�GO==�Y�=
�[��"' A��xH�5�gK�z�����Xo݈&qe_�*yi�>T�k9�*�����e����T�G�;�e�d0��#����r�Ɨ���4�������Ղ�nc�U�d�*%�c%)��(HA�§�
�����i��jms2�歎O/,~Z�q�m��ےh�yݳD�<�k���ؚ���d2���d@��9Q1���=>�\��=|�w�O�X�ٱ����c��	nd�`�_�`�֘*�yK�/�Q���b�`�[�sq��D���2�f�l�?�y�1���X@U�L{�D��U�	A�!�����̟\f���x�ߵ ���jU�=��L�VhW��e�:�E�#7՝�Hn���Ơ��BL��L�w�y�+Q�/����!M�F�1i�J���}��j��F�n���ū�I���y�D=�Q���iT�e*Ts�{��P�̖E��jL(5�
T��S�J�1��{�q�$t�p&�늏��Хnx�$M2�W2��P���O��m�w6-U@5�L*q��߳�=�a��n�@�ףF�f�D���bu��Q��ٛ��p���8�H���(0�ә�2@ý!S����L� ��^��i)D&���e���p9�E�I`�Ax�4D饐�A)>�sɸ{����O�?T���,��A���"W�0�3�te~FIOa�6��w��Sy<��Cm����Y�����J��g��7XK�sY��r��ux���#�N�)�~����;��̂�*N(��=1�c�=�hٶ9�e]��<2֧14
ÿ�R�S3�Nag�����*tj3k�~�p� ��'�a�J�ZzC��-$1m�]������.\k�{]���y�o�1ݱ�Xwk/LX�\BW��0�2*�C��Y��;.���پCsZ�&}��UK�����Q����k"�ȟ�.,����Jm��e��O)�gÇ��VS��>;K����4�\e`ӛ�����?�F�{l��k�_'e%ga� �O$Y�v�<�8�Gy��V�Aܔ�Y���F���� JM������ͣb5��}�缾�:�DyZ�<�25N���D�.d)2aI^\"��K�%�I�v �� ��P�3h�#�x��Rkٛ\2M5<���{�����ۗ�Ʊ�>����x����(G��EC(�P~��U��������58_��Tn�Ch��F��<���I%ʹ�������ڿ�%�UX���`��W��\؄i��2V�ë��+i^�(k���鸮��]���83EK�'"���?�>�M0� �X	~b�ښs��mwo���V���`�]���'���S��Z9Q����_�W�<:�]��g�Z���z�p�����6��H�H#0#Ҡ�d�E��>�\�0t%����V]��yܒ�l)�ļyF��k��)p�\D$��I<D�;U���_[���|��zM���YAȴ�2i��ju�1ry�7��ۓ�߅����Uw@�a��uN(Q�迂�#��������վ�C�[w��1EK�7_�o�c��^ɚ�w�760$�� }>7��D�����ά|�W
JV�N�1����������aX��f
?Gc��L�A���7*�bR��#��*�5�Q&p:�� ��qt��G�c�IQ@���$���jȉ+7�����N��,��b�X�X�V���،H�����|_��~q��_ǯ�����&�\so�z�J#�E����jdOl�:`����X������XJ}<�<I�����f\�Lh�+�c�d6&�@dr�g�m�cET0��I���}YN�X|��C<+@IlOR��9�Aź~���e���BD��ݕP���9/.�nL�In�d���=v�xk0^M�&Ǡ��"HnbG����U����Yձ�������� �S��mf3�j���lA�7�K�˞�M���N|�'T�!��F�/� �~��u�LW��Hp��J}��\���;��J�pϱ��a#��M��.�{���P��d�x(��"+et6��2��$��@|=!c*kPr`���u2j����������G(xY4��*t�N��! �n���t_\<�Ltk���ڱX��	٦f-���@և����2z&rX��-��=�VV7|o_PB��*w��u� q([$$���e�� �P62&:����l�(���1!��7��nq�ԯ�������n����^���4{���p�=�������@i�gdڊ��n�a����1��U9F���ie��c8ݭӲ��R��D((A>QI*cC�F��^�G��vHqQ���aQ+u���;z9�e򏖮�Jgj���A/�<�9x�iJ�@~;\7E������Q�[zҘUץ�*�j�Y��tQ��Uc���e+(>Ol3���2��"�'Rjv��<%�%�ar@�M�*<�tL�b��
��!�EE��,W��o�]r2$�4)L-�(~'vUa� @�;��h��6 ��&���U@����hχ��vn�9Q��&l|<�jg�\��Dau9'K-�d i���t��#�1��5��0"�[a�I��om�4@Qj�0����5X�5�!�'�9G_��D��U��I�+�$�}|Ջ���ٟjՒ��|�(���l&Kf�F��g*�,U�a[~����!�_W����!��.\@�oO��߼f��^INp�˥SjX����/��5T�,���S�-,/�v�{\���.z�{�lɖ ?������Z~���u�/f��u���	GɈ��CK�{Ő�F*ڦ��
�Og�A��iV��]��E����	�w��C�����p�S����t� �˵����b0�S�?%�R�ێ���ԛ�=h���v�c��pl����}�k���"�,{�s����,k��[�ʟ��,�W):+V0��;ɪ�qPD�?r~[�=�f��� ��+2W�/X�B�Sr�I��H�.�-�VZ&#�^�~��p/�x'�}�]z�X�RC����j�����F�Ns���^���۰�N�<o;��~I�ak��9�|�����k֯��1�������B��K�R4��u�%���!@t��x+v?�o�"��[����6�;�������gO���\@��&_��\;�}3/P��<0���7ʑYj�ĤU�c�@��.�E v�5n^ũ{��m����-1�]���Q3fo6'ϗIg�[�ؖ�5z�,��pn�!�7]a���%0�t ��T�*]�Q�U��}��>UK���z�ÅB�ӭO�-FR�+�*�!�'��I�[�Go���a8���.k�RP���ى]��V�Ǳv���ب8<�!�H����!���t;1a�
GY���g��:f���mc٩/�������Sw{Bfvy\���PeM�׻��.$�.p��<U���H�╼B�6��gi��}
i���i�e���{
?uv|]&d{��8h���0!7>�I7��G�^6�
�7J��3ҚF%��drml�~�|�A����h��%�u��d������gd�\�mH��K-R/�n,Nm�"��G_�6���,���/�g�vA�x&-\�k[�ɍI��V�`/�v%��\�$'�汬�/�vE�r��u�K��B���oj�*8�j�͆_F��IV��u���^E�\Zu�/�Ws�P�kIx��>�ɠ%Cٞ�uWF�r{d���I�oign��<nM<�n�E,��}#���L��\��֕��ɣ�`)�b\0=�j� �^re�Cˢp���G��Ė�������Orc�Z��|��D-HC$/���)�Xw�>W���l��7�B��`�S�Kf�i
�(ݾض��9*�����C��
�{�n�~\���=7ҚI����K��sU�_8�"������|;�<���{5����E��(�=h�����׼#!V�nj��s��:3i�0�����ڂ?nH��sL�A+5	�/���I����|��7'����ˌ�2��q�]���fl�6P�_/�j�Ͳ�S�*�\����8�E�z~�5h��	_�'쫿�nMS��?��g�t�C�׮U���[_���8,��%�cϷ���(Fco��Jx���*���e���?���<��C�gd�3�~���X��j���� ����\cwD-��V�ܠ���i��ܟ��|���,�V�������v��9CE�N:1��<�: ��t��I﷚�"��f�8$��B��{���^�0n�?ZK�Q����qvVl��@R���0o���_#\y�X? l^�����`��@�}��iʵ؃��sVus~�˵� 	"KM4W�2t��3Pd��}���pUaC�0������v��&W�a���͟U�viU�=��~`Ս	���c�޳�2߿s��W��5*�d���n���2<�Z��o_�c�R60��p]�?���r�Ӡ8�A�T�A�\prJ!ɵ�[����a��+�sA�~h�/c�&�a�Up:���=k FV�$;�e��E���T�X0��Ӡa\$�7_��qlM��F��X��y!N�V}����mA��R)|�;5�L�
�Cm�����O�ZЌ^�Bm9�3*[��v��}]v}@%���{
î_1Ş�hΔQr~��6�h%�-Sǖʩ�����Ri�����&ʔ�M����>��?��\���F=��<`�MDU<�.�m7ve�1���_���>4-~L-�L���S��v�C�!��: QbrT��JW­YE.wR����X���$�ْ�)��~��rRy�Kb�U�eL�Ñ�Դ�{w�SߴP3����^��g�$����m���O!�|%%'6Xk�OA;��}�K�lW ��̇�#��h%��v�`ooH	-����jh�"/c��?nWi#&��.���;p�4@i���yH��\�,V�����Q�Z� �K��A����ϜMҗj_F/L��3z����p�)��K��˶�y)�8⬋x:�s̿|.X���ϺL6�LAA�Zs�g���!dJ@���PA�Ä�n�A�SY���֕�`��V��ы���$�3WMw�R%k��I��ص�!6�dՆn�
ջ�HӾ���,��؇�IZ\�W��U��o��o�A+�"��`x޿{꧛��&j�@a�^o�����Ҫ���0�|���57���0�ԪKk}�.���_�{��y_��X:�Ir�Bh�0߄ՠ"��"�����S]{f�fm�X�3�P2_�5���(FB���� )��v���?�.�'kz;p������k>��u��1rzbsuf�٭XǦ؏��Ά��,a?�ť���K߭I�����@��4N���nV���M�ܹ�?���hl<�m�Uù;��p"��C�7K�L�q��Si"#�| �8���%���r��o/j"10{�#"$o��^?':2$�_;���EI�n��מ�ٌ\Mz �#2~��}��1ΫU���m'�� X4��jQ4� lb�J�"g������7h��TM��|�j��H�Nb���0x��nȜ�룊}��+V��?�n/����A?��������qՕ��g�C�~���C��v9�\��$Z6�W���68b��y�?�/�ڼq�q$@�|sƘ-_�m�Lx��&&������b6�h�fˈ������%�@^9�:1~�J~�����˰���ϛ�y��7��H��_BnkpU��25��q���R��v%�Yd�܅��;𕿵��U:ɖc�a�
Ђy���m230�)���'��M_�%5��3u}mힴ�i�(�O���q_A?�4	SdK\cT��0ȑV'D�X�j���	����L�m�j��4w yU�f�Ø�������*�_x2�5���Y�?���K����5����1ff}X�Kԉݨ�����"�^~h�������dy�P��ı2�Y�9.���=O��5_(��?�u��֡��a��"7�* �ZWΥ��(<y�)h��w����\�c;���^y%{z��R���~�$"��'���v��@�x��L�	ߚ�e!�Y;6�	�]^�����/��d+M	�n�agC��f��b�~�1-)F#Y�'s(�lY�7��F��NC�{Ny%"�B�1r�;�kJ��9g�O��2+x�c�����[�L��s��_z�gҤ��L{�y�o�2S3��i�xC���~��qoO�ݮ֡t,G���qB��kX'=����x����Y��liwׅ���R��`	F��}��ƨ�A����G'/G��\��˃����F���y��*��B�rЖ=�v1���ݚ���b�������o.M��}�đW�p��׽�K����(U9#"�6�
4
������W��d7�*�.�GF�{�d�]ʏ��A���.�1�M/�?�@6�(j�x����hb�|���1��>���*��T�!�çv��M\�Z-�����fA�@���+��ӈ����:U�W�7j�F
//(v�3�)�ϸ:��pc V}=��B�pW�cSl�`-�+^��k������W0;��V>�T*6���ٲ�,�����zjI#�v��o�,�SΆ��%Yf��L�On˥�Y5Baq���}M�P[�"r�{AU���<�	�K���z��jbV>?��[d�x�*25����I��fQ5�LԈ�6�.��x��V�E�����	ZD��G����h�L�¡l�:��/us��P�Fw{MX���+���N����B2�X���p��m��uK���j��*�yh�j1�:�	P�xIQ����x>6q���aV ��J�x-�ȉ�E�N�x�MJ�.��)pl�=�Y�� ���<��{g��of|��^2d���WWkjp%bαKP�Vz��P��$K:i{��]����Y8ކE]U൳Dgg��S\I�J�1��J$�������o�b�OS�Z�*�غ,���Z(�y��ҝo�*�v�1�ຢ'�,vs��߸���%�W��(�� ����fH}�E/����֓y����G�.]f�'��Dq~�N��=һ�7X?&��>&��JN��
��ejK<�ŗ>D#l�38#�[�_d?Ns��Q��z�`�����,{��"i��V��.2gƍ6([�͞,4h�@5�;�nL*�܍X�R������tB��(~�H@.�G>��`�֏8����|M���u��+sU8Ѧ�~�#��C֚H-HT6�]~2VAאZ�Vϗ�����=jL����2���,=cCR޸��L6k��UN�Up�;X�m��KIˊ�n���Ywb�a>��`�Ы��@�D)<2E=�3� �(t��9��8g�
m�_%�����r�����y{ ���(/)�*h��Mz�)V�Fo�`sbVfb�{G_�!��U%6�SLi������^]����\\L��"�?��IO��U�����T���XZ6ѺG�h�혽�7Z�O�a���|b����6HSh����%�������r�^��-���U
+@���7ؖE�Hі�_"p��h�gP�O�p<��/�]N)yD����Ȼ0IbTz�V��/�l�<1��7v�C#aea�� �jꁏ��q���� 0W[w�=���]�A���Q^�x�zB-J>4 �.z�Vҍ�2u|�����X���QM����K�-W��iu�8��/���Zz4�8�7�Zb�ߝ�/哌�����k��Ś�H���6�����5�� [n��\���#���T���y�~�'jf�v��?�C����Q<4�����h���;f7�2C�P7�8�o�S�`l�Uh��"O,v���X��:S�Z�5���Q.�b.$���`oI]��>��a�F���ߎc�����1���Ǡ�-{i��i��b����Q3e��ܷ�l*�*�͠�ۯ'�G��½�%��N���]EǺ�:�|׈�{�-���3/41|�!yFe^Bժ� �{�a��D���f�Z���g�����;�⼆��>y�X�c���1`I��qG���*C	���nϊz1�`Qh��[0-��0e������,���DѰ�7%o�^]���M,o� :�A�)E��]���������������F����qV�O�K!n����|K��� �74a��^�J*��(\>~��;G�ͅ�u�^�I�&���q��%JՕ!"_�4��U������V��lz��hD�	��a��Q���zaZPB�G��`ο�٥CjYdx@��{Kj��N��'=�hy�òg��[^�H���������OaK,F��Z�E.i�+-#Y:����
�'��iRLҥ[�f��z��3��@I�%	��4��h-��G�3OP�b��=`Ə�(��X�����y�a|C�G�� ��2&�?�*,B~��� .��╷%-QU�	I�fF=_��sE��wB�L&��Z����H&>?�8���N�\> )��ϻ�J1�����{�{�V�u}e[g2*$�4���z��G��A���V������nF[	.u��hv����/<�-�ٍ1��{�,��U	?���1Bq�=�l�����ۗ���'���ȧ32��f�2�BC��	E&�6!Mۏ8i!
�)!8�$��_*���#��
��-��9���=����y������Pg����k^9�DQȼ�f+x��x(u0o8�N�MuU���0�{���e�ý�R����lzI��^�T�xu#B���Ög�;]�P��F�Vɘ���OO���-����U
�����g���ԩlF-
/��Y�L^E��U�K�%Cb�A��=;�]�fR)�v��ZU����羀x�GP3���\�$PNs�ض�=��4^�
�Ȗ�#��������zv�@d�W�D�h!g�w���
�#eaL��S��լw�O���Q�6k�C͓�s�����>��@i���3m� 	����{&�t��!xk��)�<��o�Cp+�F��
� ��2��ɹ�CL��d�.���55��Փ���\�\�������^*�T9:N��]M��d��̄⒛�Q��r�;�D`���2��QN�ӝ���<�hc�Ԟ���ޭҀ��x������ڡ�/�� y��k?��K��s*kbR�.��덜��{w�WCg.!�A*�byjP[����ɪ����T�=��}`BG`ӂ�e����1��O':dKOE��5E�' /���n�S���Dt�j��FQ�[:Q�CK���*'�O�$����u����~�!gc}�5���3)[��,