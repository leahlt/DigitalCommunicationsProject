module part2 (CLOCK_50, CLOCK2_50, KEY, FPGA_I2C_SCLK, FPGA_I2C_SDAT, AUD_XCK, 
		        AUD_DACLRCK, AUD_ADCLRCK, AUD_BCLK, AUD_ADCDAT, AUD_DACDAT);

	input CLOCK_50, CLOCK2_50;
	input [0:0] KEY;
	// I2C Audio/Video config interface
	output FPGA_I2C_SCLK;
	inout FPGA_I2C_SDAT;
	// Audio CODEC
	output AUD_XCK;
	input AUD_DACLRCK, AUD_ADCLRCK, AUD_BCLK;
	input AUD_ADCDAT;
	output AUD_DACDAT;
	
	// Local wires.
	wire read_ready, write_ready, read, write;
	wire signed [23:0] readdata_left, readdata_right;
	wire signed [23:0] writedata_left, writedata_right;
	wire reset = ~KEY[0];

	/////////////////////////////////
	// My Code
	/////////////////////////////////
	
	//Required helper modules and files: GenericModules.v (VariableFlipFlop, VariableDivider, adder) and FIR_filter.v
	
	
	wire signed [23:0] filtered_left, filtered_right, noise, noise_left, noise_right;
	
	
	//noise_generator L(CLOCK_50, write_ready, noise);
	//assign noise_right = readdata_right+noise;
	//assign noise_left = readdata_left+noise;
	
	
	assign filtered_left = (write_ready) ? readdata_left:24'b0;
	assign filtered_right = (write_ready) ? readdata_right:24'b0; //Transfer data from read to write when ready_ready is high
	assign read = read_ready;
	assign write = write_ready; //write input flags to output flags
	
	FIRfilter left(filtered_left, CLOCK_50, writedata_left);
	FIRfilter right(filtered_right, CLOCK_50, writedata_right); //instantiate filter modules
	

	
/////////////////////////////////////////////////////////////////////////////////
// Audio CODEC interface. 
//
// The interface consists of the following wires:
// read_ready, write_ready - CODEC ready for read/write operation 
// readdata_left, readdata_right - left and right channel data from the CODEC
// read - send data from the CODEC (both channels)
// writedata_left, writedata_right - left and right channel data to the CODEC
// write - send data to the CODEC (both channels)
// AUD_* - should connect to top-level entity I/O of the same name.
//         These signals go directly to the Audio CODEC
// I2C_* - should connect to top-level entity I/O of the same name.
//         These signals go directly to the Audio/Video Config module
/////////////////////////////////////////////////////////////////////////////////
	clock_generator my_clock_gen(
		// inputs
		CLOCK2_50,
		reset,

		// outputs
		AUD_XCK
	);

	audio_and_video_config cfg(
		// Inputs
		CLOCK_50,
		reset,

		// Bidirectionals
		FPGA_I2C_SDAT,
		FPGA_I2C_SCLK
	);

	audio_codec codec(
		// Inputs
		CLOCK_50,
		reset,

		read,	write,
		writedata_left, writedata_right,

		AUD_ADCDAT,

		// Bidirectionals
		AUD_BCLK,
		AUD_ADCLRCK,
		AUD_DACLRCK,

		// Outputs
		read_ready, write_ready,
		readdata_left, readdata_right,
		AUD_DACDAT
	);

endmodule


module noise_generator (clk, enable, Q);
input clk, enable;
output [23:0] Q;
reg [2:0] counter;
always@(posedge clk)
	if (enable)
		counter = counter + 1'b1;
assign Q = {{10{counter[2]}}, counter, 11'd0};

endmodule


