��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P����z��{}H���_Q�hФ���]xy�0�|s��9߼L���حe=�3�����Uh=8G%�t���n�4��D�cm��zۜq�a��?w}HC�#u¨�`�L�Cަg
WS�1f�k��Z�WЁ��ehg�+ݖ��F�	Y���җ��2)W��Á$��%��-�B���C|;\�z�8����P�����`��:���\���c��E�14�QC4��l���&�d�2]JQOmF����q�my%�!��Y(F�v騜���b/�a�s�c98�o0t�w����M�Фk���3��u������tXv�8���$�N�垐l���������� ���4�?}#�+HMعM�49M�����&#�C���?*w<�SQR�XTn�61qK�M	�{	t�u�Q+�E���8FBI ��j�m�U�h��_�rt�3�!�׈/���"�#�[�BO�#pϐ�+�I�?O8�P�g��+��~�5�W���蹋��oС'� ��Ag��j8�
���QF�����^P�K�Ңå=pƹ�a��I��!�oýN�C�սU͠�+��P����T>�_X �aۉS�uU����3ԉ�s\] �PHQN3"�a�͂<p��nM���{T��'��_�����t嚿���
�_���\q�͠~��@��Pm�`�����OQ��8	��Ռ�\�h9�Q�
��v��ZV�_<G�J���~�,18�h�h�r7���0n|�Pꌚ�r�LG'(EwO��j���:��847������ۯ}x��|'��'��m|��E���`BO9��C�)ù��f�����M)�>}2��3���K8h�� '� y�b����������b*�Rq� lH�"������g�8��!>�KF1t�}�s�x�/(|��>Cr������߫��&.��ȧ\�� tGv6栠��[��(��6�S��#��:_愭t6ߛ��YZ�
I.&�1��Jkt�>#r;�>z�18Ŕ��Ơ�����Lu��T}g0��1����&9��J�3tn�bD!�/@$ ]�������l�a5�����,�bҮ����䪴��JS'-�4#�ʒDqcR�S���0�\Q~���t,N2�d|��n���=�%TC� �ީ�ʣ?ޛ�$c;Xu~��U�jNWA��/k���j�9L��=�o�����DS �	��ӊ$�Є؛�֊�cx�F.8���1t��af��a���v�t]��^��`�<� ��U�Vݸ�S�œ:dy*w�p�Km���_A�b���P�a/7-��=p1
��7O~q�q�d��\��;8�CVi��f�Ba�\�m#������Κ�ٽ"� 7�}Z|�1����n�BQ��0�nԅ�5��!�O���>Z2L=�h��q�N�^b��Xɖ�3DI�ܶ�0�c��S����P46�g��*�V$�����1G����&Mb�8S`fʩh��m4]��L!��8��,�85�/�B��%��FL�8R/�b����f��l5���bi�HOҽ�gp;�42�tiZ���2�8�;Q>�^	�^���s/2��V���E�:b�C��bls�s]�((����D0l��0/�@kE	I���z���%_��.������[O#�>4`PWH�p�ԿT'��b��U�v��������Eal�[X��el}	�}����Hn��J�d��r,2i;�b��1��PWm|r��h�a�>�)V��������d��Xe�~����1
�f$�^�� ��x�ˡ6��5�	Ҁ`4$��^x��Q����F��B~{�����
95�-RAoe/��T�1��ͯ�(�
��-�$��;�����(V���g�m�����<n����`Uj�~QxX=�iUC�.)�~KM��Ǵ�9���ዑ��<1/�� /�+1p�C��%���Oo86��#yb�e&aFΟ�"a�H�z=�����}��{��8M�V�sy�"��uѡ��{�Q闦��BȀeR��q�Pu��S����Eb	��B�J_h�7v�('��n�Y'��?/;��wk��KvY��=����^8�<#���Q����Cv��^�S�Y�Ĩ��K�({����������}2�7�t��pP�w����N�uM���(y����1�aK�5;�g�M�<;ٙX=�nV(7]�7}�U��z@���+��8����T���j��N�!tcf#3a��M��Ƴ���q19���|!|`o]v5�d�X�f�}L����s�����߬Jt�4�D\q���a(U�i��ST4±=z��b�ض��h�����Z�:����S�����Z:nj��,����B��S��S�D�6T��Dm&o${G�N��mh;�!#���/�V�v��a��}�WM���C����Z�=�5�����8�Exx��;�{�
��!�X`:��Q�RͿ�,CB�NiX�����	�b> �������B@f��m��a|�(`�匈��9sS���y��1���烳��#5��3w+�%��~rE@��6����b.R�L�]*����@�]��d���/�aro��̴YNy��`��[j	7�T6�S@�Ke�	*F0$�KtVP�֥��x f�K�k������<���Hc�^�K
+$5�o?�<O�D}[�'���� a� g��q*PD�c�[(��� H��n"��7��I:Ҋ5��I�*Օ�|�~�zR�O�.��Y��t�T�[x��J衽�r?(���H������b��&�����Q,Ti�D.-�k�~�nZ�B�] y��;��
^V�!���g(.=@1�?+;jrG��Hh��\ڱ�j��:��	�wk+}E*Zuf�鵉`sE�Z �}��Q~��[tW�n