��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`uW����=5���2�k��]�~f�R�O{�#>rv'5\m��P���k�BL8zwg��+��6>��!��=5��R]�/����G��r�4�	�@�A�GT"jH�ki5�1�Z���h��Wa�A,���g��[
&mF&��Գ�Y�.!��� ��ާ%��n�|�>�j��ؔ(��[ �)SRs=C"V	
l H��/H�kfa�q�~%|���-s�y�<�w h�:}�+��CM���T��V0?���bv�jnD9&W��U�9�4�t��� �˻+�9xv�;A\�#�;r��@��A9g_s�6-�������"w�z������8��r@���;`\��ٔ�m�jZ���|Uh"z��9��$��Ui��c��M�jſ��[��r!�b:�����gRa�Д%p������]B^���T�z蒻��qV�J��O�h�rs�S�e��QIP8����>�� �k�պ�e~�B
�͜p�O�.�g��f�Jş��	ox��U��b��@@�7	�M���Ir�?2��d0f�үy��"6o�,[v�':�*_���a�1��r��y�9�,�t@�8tt�_�R�-,stVxYui�Y�����8A��]�6�����MBh���"J��8�t���^�.��'���)~�	��T��8�o�v���i^F�hr��~&J�^��ͳ{~�߰шe"С��)9��D���Q<V��uf�x�K�X#��`��ߦ>�e�
Cz�{Q��<�%��F�y��&�SÁ N�^�ZX�\����/j��<e��]��8�ᙚ����]������;��yj	�s`��R��y�I˦qGI�y�O�U�u��� �_f?�?ٺr�Ҫ���'7��4�r��<H���;�{��e{t�	������<C��V�gh����05:��d�[��W-�������&:#VA�L�z
�_��[��u���b�����t���q���hK)� �l�(��PI�X
�ש0����h�kѧmm��
���4j��1��V{<�N��I��`��}z�ۙ*zK#-u���4O��[�
�R��-�+���V���P�?�N_҈�@�F��NDeX}zu=,y�&6Ƭ������˸Ϻ�e�t�{?� ����G\�+.��g᏶��S`L}���?�N�L0��������f�X��@�9}����#��Ch?���mw5��ٖ6��e�!���~��+2&�@��h�x�7Q6�e)�G�F�,�Թw�q��lN<ãS�wE���Ԧ~ΐ��L����hj�y���)�y�j�4�Np�,y6԰����N�B�[�mk�O E���(�/{�3�f�i~w�ڭ]�2�4\��{X,�#���<����w��L�o"��� ����PbSĆm>��F{����S4pe >\FX]"�(<��X����Oٌ���}�z�ۚ�ڏ�,qP]9��(\rB]YV�)���N~���\}��7}�M*�Y�[/�I��~9֚{�ݻ�{�^���*�_���ӝ�����q=;���Yۛ����HJ���!z�(�U>CX|��+:
q�\	c�H��f�t�I$P{��B�Ϩ�lf��U�w9*�oԮ�{���oa]E=gO��}\����r>�fj�����89E��VfB6o��V˭����i<��IBvo83�zj �6EoT?@'�!;���GR�Lx��h/^J�{N�0�t$�7�-��&7x:��m�Қ!l�Lc�ݴi��] k��̞�R�}� �m�jy�o��o�!�>�t�A���@Ev4iP0���.>�2��[��Z!�adP�(
���w�j=U��+9�Ӹ��hs(�(��v)�?��e/Z2���<��`ܠ*��L�)��Y�_(:���s=y?:g��5�8Zs�%��D�K��&��D�hc�0ĊT.��(IK��]��P�'Y3�X�� �����\�!����
ע$�����"l&Ģ�rSǣb����E�1�&l����8�2���4�1qjzgE�>GW���*�+�Na[���a񸋤[2�BcP��.)z�J������u�H}�6���\�p'�t,ѝ~ "F�T��~�P{Y���b��\�� ��r��Ô��ε�h���v����wT(L�o���P�c��꒟�MN�<@��N�^��@H����IjC���x{�1���H��-/��5�}�?��c��qZ��z�-���o0�ɼJr
�1��_~��D;=�����{w�:ك���)���\;��IKs�;�%8�7�2<�jT+�*ÍH�g��9�?�{��&�MSm��"uE�BH���I�S�8��P$i@D��=��C\�Wt��<i�4��J�����]�-���޸I1��J����!;O�av���L\NC�V��*��E'�2���y�Peг^o[�SY
�Þ���x��y�Ȋ�劊ǿ}��?�E_C�[P�,�]g�b�_&���_��DpoR/�!p�s�@V!��0���0�Q�u��kr�>`^_���3<�SPtԡHʨ#p�s�Y�2x�Qu���|���_�z	�,���h��4V} t�rӤ@��xy�M����ecr!R�=e����j~^��tVc�> �^�G���h)����MVQ)�iHι�v�|�>|�sM����C���P�|GIUǠ���˺�f^�r����,24?9����I�W�~�|�"`��"`)���.�m�R�ߡ�f�?�.vN<v�;p��[/��-�8�š�������`kC�±&!b=N��!G#=��~���2�Z��6{LL�n.�Q��[;ʡ�����|s�d���=���{%���6�#�2T�F��D�
|L��An�r�o�x�tW��iҷ�#)yf\�����Һ\1����-)�^x0�u���LH�Z��r�/�n��͡�Y9э�~E���M��æUD���k�ʜ{lJ٩&]�)���i���2ӎ`�q��M�J��, K���� ����6 �Lo�	6FX�9�E%7�u� ��Ф#�_�T����#�o� 
���x��k�ट�l2��Õ:0��D	�J�"��X��vYg��D�W��+��Т�����q�CO����D�$�F8$�����h:]�ěN��T���5�ӳ
�,�g&����q����^������0< �)|#o|�!7�A��jj��İ���i饧�������y�ۚtk������d�W!�wtT�,Aq��9���~]�=����m��LXW�A)Sï�>�ޥ
,�F߯E*̫�I�Ɯ ��.�դJ-��phP�p�C�.d��y�t(�� ���{9�G������!��V��D�k�m�*=�����e���3�r�����D����Lw]L0�B^V#�5r���պ���� ��`�:�=���'˦qBU��0���}�B��s/���I�lJN��z��j�Cy�w�-=��nF"Pˇ$G~�M}�&%'�������8$��"{ۇ�V@A3ŢƗ�D��|9��g�m�mʡ�Ҩ���b/�Xa��YE����p�M��ŝ;��!��֤,V>N�M�[q����r&�/Wg�� �zo�A�/�1��Loڕ�2I-��TЩ�6����/���T��@n��Ѻ��e],�_]���"�_�l����\���F��c}�l����Ǫ���V��E̓%�vϡ�̱��J�p�/�������
�� ﰌ�L�r��1��3�)���@��4F:�9�L�!�S��-��J�Z;��.>�f
ʅ��U��Z�ɮv*�+�W���|6�AVkA[J�-N��w0��_��}�Q˗.��.]�.u�W�JW�#���ugzHDf�����i?���^H�m���
�]���Y5�|�Z#�����z���"B���f�+����)��1�KSݥ��ͺy��m���Y	��3T�@�Q���KR���=����Qr ���`RCk�J�.���6���}�	�.�������4�w����a�]Y6d2D��ʭ�"�@���o��C�$>���b��󎻭�D���P߂(�Rٲ��Z4\��@��'u�Ga�/�T-:螖t4 ������h*���2cu)HR�5�ܧ�yWS>��t�J��:���������Zz�F[׸�]�������>hs���=^�����y�����N�fK>��H�%�bl!�M=�\�D�r�bd��W<q�Ċ��	�p��vJ����P�������e@�$�XJ,��-D/̋6��r�r�S@v�_���U؆0GfU�G\�N�#i�~�SE�@rj�N���g�����j���䜬U����ۨ���l0�"�O�w� z8�{��*���
��t )ŧܖ���ny�ԇ:�/�W�W����9�����x(&Yd�Wn�K=A�D�Tb|)v����qL�,���Rs@L���*6=�du��+�}�_���°n��{��t(q�X�����C%{�[P��U� d-e�kY��@��f+ E��\����;{#�5�-茳 1�!yP�X1����ʀ=lD;����k5�xpr��G���l�o��;|-�2�)���f�7�k��Z����N<��	;0i{n����VI��ƞE��1Ifh�]/�����p}o�q>�E㤶%q����2f1"�퀝Wn�}�R2�5�\��|�5������E�c��[�(ڄ���Ȭ]��у[2�9�}Y��*��ﺰ����q�^8���5�� /F��.�x軦�ٚ�� IE���~Ϧ�^Z�t�l.F�ٸ��e��¸�h��%�*IrR��W}xn��Iv/cfGp�!:O�X�XΖ���j��]��P�S����EG�mU�$���D:eޖoڡ�^�\8��j�woA�@��#%�4�S��Pߵ��ܝ;�s��m}���sw�U��E �v��-�^e�������l�����Cg}��]LQ9�E�n/���%��B�����[�[�>��B�h (Y��0�L�,e�^�:�⅂�֙G�`v�e��g�K��R����,L�g)�g<v���l�Z�t���J�,�w�#�7S����������/a,j�����& I�̺�,:)a����]� ������lZ9P�q2%��:l=fG_���7<�TOF��Fʎ�
��\�'k�.�.k�^����G��~��h#֪��H}���2���Y����������fY@Լ��ƀ�,��b�b�S�Π�|�L�9��?��A=/�����09hi]!"]�O6-i=���ۉ�v���Q�������#�t\��%��X5�lk�u��S�B>�� ve��0+p��ǐ�Ju��̥�ɅN� �]63��:�0�y-����t[u�
>s#�]S���M(�>����ax��2g�D��,[yRW�Z�?�A�^k�����7���� d��8^�� �{ym}���8�t�rk� 2ɦB�0�Kb�;(>:�	�@�}'f��!���h��S��ж�4Q�rU��Ե�%���Q3B����%E����y�"�S�ԭZG�{�`ޱp�V��&����Lx=��hcޡ:�*�|,�4*5���x��hlo+��������D\�ȶ��H