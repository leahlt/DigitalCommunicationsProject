��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P����z��{}H���_Q�hФ���]xy�0�|s��9߼L���حe=�3�����Uh=8G%�t���n�4��D�cm��zۜq�a��?w}HC�#u¨�`�L�Cަg
WS�1f�k��Z�WЁ��ehg�+ݖ��F�	Y���җ��2)W��Á$��%��-�B���C|;\�z�8����P�����`��:���\���c��E�14�QC4��l���&�d�2]JQOmF2FVc/K���)œq�TS��f��7.�f_j���M"�U����� v*�����%�I�bI�������e�>�S��"l\��G꾇Kv��u|�� �vuXР��UO�6sUR�o=�B:�dw�I_�ʬ��@�^���~T�ti��+���Á`n������L��i�f��6�cu�/���t���o��<m��|{�J%�w���lErkR�{�T.����j��I_���{!o����F3���:��5��Oӧ�������w���)� ��T��IT��clu���{̔���)�ȃ�s���M\���$�u�0�����?o;q��� �ߴƣ'��$;�m�rO�K�C��+Ln�ִ��9�T>]������s�F2��7��lQ̞Lb{2�}axj ���Gq��.�~w���6{@ rny�t��*������G������i�
i|��L[N*ʘ>�\��5[��G�|��⒦�Q�,�����?6�"nj`�0�_;��TRT���}�-�ꥋ�ʹ=���:A���P���Ұ��*�XN�\NF�+����{;FJD5�eA�7�e� ܭ��_%� �&��_EGΫG�z�UBN�����ǣ%r"҆*2G�����F�î4���?N�&���#�B����4�ĘSI�dp�n$ם����K�߲A 
/0}z�H����=�H�^
nMݦ�|�̼[B�1f�<�[a�/?G^�����fi�mϱ{��~�(av��6o���汿������jTJ���τ1v)����٭P�i����q�6�,ęLW�I�p�)�����m&,���H*��3+g��MM�����
�F��q��&��h?�t8�y ��Lϐ Aj����Tϼ�+ZV�IKy��X�s�j�)��;e��4⊗�,�e1<w`�<]�[Z�3�ITj�OR�Oܽ�ߖ@��W��'j�ͮ/�����[XsE?+ʴ;q��o�J0Ӳ��\mr��6S4���g����}���7��/Fr�H� e@)d)���}S?{�˖g�_�%��*���A�Cc�׼(1���%V*O��
�n ���n�!;'@ݮ�}��w��˝�Z��z�� �m����KA��������