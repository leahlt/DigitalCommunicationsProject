��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P�|5js�[`F�q�t�(���(-jp��
�����-V�N?�;�� S���H7L���S�w�Wj�K�DP2�_K�=@�%��՜5�A���hD}�ϾSlI��iͮ%��h��Ԣ�^g� �lT���A�����}��LY������&�ւ#�aZ�p~�J�YGO��ra�w �_7o\���|�P�;�I8��ѣ��Y�b.'� �yh�b#�������To�{��`˄R�K)��2�Ah*��U0��<���75'��h�B�-�z�d�̮�۱�T}�?�K���ӹA���&�"�bt	]~��/���^[�;���PݴQ�$
�Z��z��&Š��s��>-��,�U_V���m�D�����0�	�L
uۻ��t�5%*���4pg�:�q���f�)�4s��ޙ���Y��Q�����{�z6����*΀P�	���f�C
T�P�ݣ@K�~8�Q�2�)eчmz��N���
��� P1X/�����̃�8��|�{�-��qa#^ۺ�g�_mӄ\�(��̋����֞��l��4��G�<<X���;�����bls�����i��)���A��bM6�]��N�O��ERz�����˘}[�¯Oh��|!
B�G�Dm��G��1occa$�r��w�PT��MꝘ��dW=���Ho����m
�]]*��;��\��D�0nJd��E��|�&`���;5���B��"����F��0�}*|z�&�m"���D�Č�|#.�cG���0F�������U����[��8����[wP6N�`m/}O�>�㛞�������r�!���a��s�T��n�+B��v����#y��0O�`tF.1�G}��϶���W��$�tDx�85Ĉk�ĉ� �܃[��NO7EB�iY�d5�#sD��(-�:AW��1C`�,)��Ŕ��b���
lE+M5�E�T�η�I�)a����W�է�
1H�<�E:^�P��`?�42B1�\���������{�4����y����A�>Om�[Z���� ���!Ĉ��X������	}������В� �cU��a��(�:��{�A��]���i�m(���k~�s�} ZD���	�d�q�Z�%F<�ߩ_��s0�,Q�Z�~�M��ʼSZH�H���Ъ^O�é,�Za^��K!puHf7^vD�u$�h�2��j|�
�;�ڈ�n�Ƈ�Bj�'u�5�pQ���	��j�cMQ������y�u��a�3k`�4`+��'�ۦi�5tt`��@�z�B٣�9��@T��E��W��:�r��\1�cq�s����&ڞ3"{_H�I�%���Ƹ���ci3����j�֡(}�
�@&�P�b8�E�y�����njM�[cU��߹SeA�
����h�'��mƆ�Li�I�a����w9e�
i�g#y�+��PY���KzE� ��D����Q��������_�-�W�jsAOE���jKV����Ε��;��o�N�<!���{�_p���ɇM�;��YN������)7IX��.I�pMJ�ຘ���ˑ��V�JM�v	�ؕ�'��ǝ���},�G�9�|�I���,�_��Eo[�6�D}�Gq���3xiN�WI(96�z��^��c�ٰ�'G�W*�>�b9��0�EUI�~�G9�1�UN��&P2_�����?���1�s��A$���k:*cT��� ���v�!.�t�L��7��c32��L�1dZ`�T�Sg�
�)�Ѣ7W!������Y�� H �˲v̬|9(��bDY�y���~q�Q���32r���S[c�TU�q�V��=�бq`�ԀJ����]U��zL���aI�:m������$G1���ër hn(����oO��=�W�t�����ԘI�P���Zm�~���z4`='w��>� V��C�a���槻n2&�	�͟$�B��.m5Z�C��t�[�^��9" �5M<n���>uf��m �c;yb��;\�aZ&������ȓ#���g�9��D��l��bJt1:�q�=-��� ����I�$�Ŭp��>�t������-g���G3��q�n�j��P���%���!�O�`�c�A��d	M�����_ʣi��3�AZ�	»����ȯu�J���x�)a��M���Ӈq��/v�> Y���D��2D+�њ�l�]����9��m�<����2ª�$��/��Lԗp�hX,7	���VZ=�P�V׌� ȘI3T[��ė{R�޹����C��\��g��2:�6Q2B2��*sa�������#�h������!' ֱ�Ɩ�6�i-F�J��=&/�
h��D.�V�ݣ�)vX��2��Ѹ�<�C�(��k ��CR9k=��t�S1�$�C���hn����D[mWo;�uiZ����0&��g����c���7�Fv����&�,P~�
 ��2]~H�u�"��6��m	,r7�?�p��L�"�dS$��^a�7Gˣ�!�I	�֨���G���رR~|�&ԡՠ���fBF{�3Sv+߁l���
w���K�E��>]�� vl?�F���I}�m��h�&@v���z*e���=ޠ���ŉ�]�ŋf�)�Y�֪Lɠ�R>4�%�z���16��#�*��C錇�
�0�bh�2��\�yY6d/Gގ�L��l�I�O�٨[/��y[L�oء��-_F����7b��@a碑�!��:^d�{-��L��}%Q7�Kv�f�)���:�rT�ꄭ5�E���Y�"Z|@��%��km��8Ѹ�d����^����:44d�TXU��aľ�D�`�Xс�Ds��9L��b� U��v���C���C8���{�'Ɓ��
*4W�V2k���>ͻI�;�����'�Fpݸ�(�R���45�f}?S�+-�咟Ԛ��H[#��*�s�DHq�Y��
z�+�c%�9�����y�{��U"X�Dg5�Pi�w��-2����鸩�yС^���\���ʽ��u��Um�-p�^���t�k+O�o�����8W���'�2
�ߒ1⾒�E��1D��AH_����-9i���;�y���)&B׻��A��7_ʤ��ά\��b�*�J9�ۜ���X^u�&n�'HK��X�M�:���>%��KT��QcN����Sb�n�V�m��Sql�;��{��y�e�z�4�����#q1�`a\}�ƨ!��=Z�M2�쩔o+���,fH�7<�^�S�w��V��ߙl�)/�%�"8j�g�Ǿ�η/�m?15��$"~���^&��m���̢��ω��
�wD�Z�*��!�5�F;_Ώ�>E�*�D��M���XC�KW�N�o!�8�0V{"����L�n @�-�9�D.���.u��_^'�����^�y�;0��׿UW�#e�\�o��%y钕��-�@�Z:����!2���8'��V�2x0����58b�]�s��3��p��}�ZO0��Q\d�M�מW�8��勉r��}��c�	���.?e����/!�h�� ȕR儭������J����tVi�&�7lY!F��tQ��A�;WO�����u�ӛ���s�4Nx踯\����J\s���B_�$[G\�75���t9d�c�����r���`��gh����JFt�;��ϻ"�cg��^���c���������r&A�V�����Ø��b��������[D:et��6�p%Be?l����3+�u������ihl&kSٍ�8��h�y}��ף�a
��uq\)�!��c9%��ȏBh �� fN$2�x?�:Jq��#l(FY�@��8h'k�J"�\C���* �"�!4�wci����[�V��k܅|oI�@�5�A��*���F��o*�J�$-�ڙ�����6�w�X6�ǔ�g�m�N��]>�X��d��'÷�������vg��đ��u9FJ��+���S>k���v�Ŀ��k���6[N@�_,��