library ieee;
use ieee.std_logic_1164.all;

package bch_enc_package is

constant CODE_LENGTH_N    : natural := 244;
constant MESSAGE_LENGTH_K : natural := 168;
constant PARITY_LENGTH    : natural := 76;
constant DATA_WIDTH       : natural := 24;

constant POLY_COEF : std_logic_vector(PARITY_LENGTH downto 0) := "10010110010100111001000111001111011100000100011010100001110011000000100101101";
type lfsr_coef_type is array (0 to DATA_WIDTH, PARITY_LENGTH downto 1) of std_logic;
type lfsr_input_coef_type is array (0 to DATA_WIDTH, DATA_WIDTH - 1 downto 0) of std_logic;

constant LFSR_COEF : lfsr_coef_type := (
                                        "1011010010000001100111000010101100010000011101111001110001001110010100110100",
                                        "0101101001000000110011100001010110001000001110111100111000100111001010011010",
                                        "0010110100100000011001110000101011000100000111011110011100010011100101001101",
                                        "1010001000010001101011111010111001110010011110010110111111000111100110010010",
                                        "0101000100001000110101111101011100111001001111001011011111100011110011001001",
                                        "1001110000000101111101111100000010001100111010011100011110111111101101010000",
                                        "0100111000000010111110111110000001000110011101001110001111011111110110101000",
                                        "0010011100000001011111011111000000100011001110100111000111101111111011010100",
                                        "0001001110000000101111101111100000010001100111010011100011110111111101101010",
                                        "0000100111000000010111110111110000001000110011101001110001111011111110110101",
                                        "1011000001100001101100111001010100010100000100001101001001110011101011101110",
                                        "0101100000110000110110011100101010001010000010000110100100111001110101110111",
                                        "1001100010011001111100001100111001010101011100111010100011010010101110001111",
                                        "1111100011001101011001000100110000111010110011100100100000100111000011110011",
                                        "1100100011100111001011100000110100001101000100001011100001011101110101001101",
                                        "1101000011110010000010110010110110010110111111111100000001100000101110010010",
                                        "0110100001111001000001011001011011001011011111111110000000110000010111001001",
                                        "1000000010111101000111101110000001110101110010000110110001010110011111010000",
                                        "0100000001011110100011110111000000111010111001000011011000101011001111101000",
                                        "0010000000101111010001111011100000011101011100100001101100010101100111110100",
                                        "0001000000010111101000111101110000001110101110010000110110001010110011111010",
                                        "0000100000001011110100011110111000000111010111001000011011000101011001111101",
                                        "1011000010000100011101001101110000010011110110011101111100101100111000001010",
                                        "0101100001000010001110100110111000001001111011001110111110010110011100000101",
                                        "0101100001000010001110100110111000001001111011001110111110010110011100000101");

constant LFSR_INPUT_COEF : lfsr_input_coef_type := (
                                        "000000000000000000000000",
                                        "000000000000000000000000",
                                        "000000000000000000000000",
                                        "000000000000000000000001",
                                        "000000000000000000000010",
                                        "000000000000000000000101",
                                        "000000000000000000001010",
                                        "000000000000000000010100",
                                        "000000000000000000101000",
                                        "000000000000000001010000",
                                        "000000000000000010100001",
                                        "000000000000000101000010",
                                        "000000000000001010000101",
                                        "000000000000010100001011",
                                        "000000000000101000010111",
                                        "000000000001010000101111",
                                        "000000000010100001011110",
                                        "000000000101000010111101",
                                        "000000001010000101111010",
                                        "000000010100001011110100",
                                        "000000101000010111101000",
                                        "000001010000101111010000",
                                        "000010100001011110100001",
                                        "000101000010111101000010",
                                        "000101000010111101000010");

constant LFSR_OUTPUT_COEF : lfsr_input_coef_type := (
                                        "000000000000000000000000",
                                        "000000000000000000000000",
                                        "000000000000000000000000",
                                        "000000000000000000000001",
                                        "000000000000000000000010",
                                        "000000000000000000000101",
                                        "000000000000000000001011",
                                        "000000000000000000010110",
                                        "000000000000000000101100",
                                        "000000000000000001011001",
                                        "000000000000000010110010",
                                        "000000000000000101100101",
                                        "000000000000001011001010",
                                        "000000000000010110010100",
                                        "000000000000101100101001",
                                        "000000000001011001010011",
                                        "000000000010110010100111",
                                        "000000000101100101001110",
                                        "000000001011001010011100",
                                        "000000010110010100111001",
                                        "000000101100101001110010",
                                        "000001011001010011100100",
                                        "000010110010100111001000",
                                        "000101100101001110010001",
                                        "000101100101001110010001");

FUNCTION log2_function (constant in_data : positive) return natural;

end bch_enc_package;

package body bch_enc_package is

  -- log2 function
  FUNCTION log2_function
  (constant in_data : positive)
  return natural IS
    variable temp    : integer := in_data;
    variable ret_val : integer := 0;
  begin 

    while temp > 1 loop
      ret_val := ret_val + 1;
      temp    := temp / 2;
    end loop;

    return ret_val;
  END log2_function;

end bch_enc_package;
