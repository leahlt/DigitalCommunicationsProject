��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P�|5js�[`F�q�t�(���(-jp��
�����-V�N?�;�� S���H7L���S�w�Wj�K�DP2�_K�����htdo� ni ��?��$";������$�
��L�I�N��$:u�|�H���Y�ӗ5��!�����ǉ�Z�il_Z�^F���XO9���D��w{f1>�сF�?�`���k��`���tS�ء9��%��	p��� P�Ő��~�oN��2��隟f d��tl$�i<�O�����_�Oh=�������c����W8�'z9�?˥�;Ff�o憭yr�n���.���#���2�D�q���%���U��K�Q�!�|�8Z�����~X ѐ.�*�N�jSQ'����� ����w��q*�Y�y`�+�o
|/ܞ�
O���&i9���ȫA;d�G�'��U�������z͛��ܡ�x5II��o�/Q[����u5)5���Ȱ1�Qdc��-y����X��edQR��,#����J�Q�����~�������Xu��ǡ(Z�D�( 0�Swy�������������\��@řd�e��-��~,��5� ��魙��z,�����}=�݀[�[M��޳*ND�k�.&�;�K��,  ��+[���M��� ">T<I�d�+~���v�"��p��ߟS�<�j����\��|��a����y;����Ei�g${g��A	��|Fƌ�����G��Qj޻��LS
_0��v��v@z�h��>�{� 謝w�4�c��^�-��k)7�ڔ�,h[��l*0��.�0�~�Q���j��7�ģ!c����Q�՘�x�3�Z��W�l���?>V�ޒw�_ҙ_�6g�+�>&�^�� �eL2����xt�i����Y�Ӿ���QԼ�MҞu�;��u4݌e6_�20;U
�n�Z�R�{����p�SÏ�x�CL&��3�j��}�ĉ��	�Ec봭d���|�&��/n��GSϻ@���ܭ��0��E8bl������k��2H�9k$�5�J3QX�翤�{$q�=�U	�������n�,�N*I�O�r�7�*g���Rz�h\�Ђ�J`�P5b�;I�'17!��՝�3�5�]�2�j���v���=���8�ls�s�H������3�}4�|m�$)�J�ú8����h3UIQm~�4���]��(��dMv��ʈq�m��W�wꩼ��X���C$��;<�$���εcS�)�w�4a:O7\���mX�_�Wvc��(�R��>E��~<���W/��D�RF��3
�Dh� �5W:��7�z�*���n�I|�)��n��NkB��yY�K,5wڻ���/+'�>-#w Ť/DS�n�*��2:������͇�=��5�r'�3S�ٓ��V� 
p2�VU�3|^��x822�C�W��S�V��b�K���9�C� ����#8-�P������C�\r	�ǂϦ=~}t�����FO�������MI�à�-��|�jX����������U�K(<P.�Y� _9d����M,@��<S�:�5Ҩ�O�$��W;*�&�ݎM
ز^�8�0�x��34�����w�=�]�mܶd��1˪�,���rK����O� f1yI�UU�B���}�� m_fS�D�7�ăn-H�Bg����7??�!hT/e�[��o9��6*5p_�oW�u�N���2j�{�t��x��y�X$?a�!a�O
�p�YAH�HN�8��!E�3��F��Ԃ�k(��&�aB���٩���޾�u`�.I;��_�D���*Vj��Q�@�@�*u]?�7����h�bdV���JZeLa���w���Z���� �2�Ţ�>uAn>B�L�=���x��	J������uR[:�4�.�M�)��\������=����� ���WA{b������銇"MK����oɘ��4��d��S���zSz؀y}`���4��������l�w'5|�}��ץ���p�G��OP�d��D	��G���8}�f�2s�X�.LX1�o>��} ��R	�`���6I`�yo]��a����!w��-���� &��b,��GȄ}���[6Q�u���{=��;���?�����w�xS�\셁�������S�|Ք����Y�M��*
�d+^�=5U��8,�|�D��Ɵ|�'2��O�TAl�#x@*���?���Wޘ��W��9��c�l1��Nnx Ra����O%�z,G�V\���� N"�F�z�r�#	��\�6�\Y�!�u�W|�@�R�L������|H��P� :!d:R�8�/e��/�3��Nf�`�V�F�"b�f|�2��H��
e�k�*D%w~>ˏ�?+ף�y�~yP���>�J�|��b壮|٢.��a�]�Z��oa����Ѻ�� �����@�]�¾c��R��}DQ�y8���H�ŉ��Y0����H��Ubg�;��Z��\���qw>��ڗ��ydG�� ��r�;��O�U���q��Ln������\?Ԕ�hY��d[�/�[x�_ѺU����+�o��-x�f)]�&���u��s�+���i��cp�d������"y?1���պ��.��,y�xWz˜��s�c5��J���������D�c�j����m�v���!����c�OcuX�̷��3��/��d��mZ��qe�H�晡<B�(m��%�:0�	�8���.�R���%�n�>��k�Գ�5��;A���-Y 	m�T���C~ڎ�D9h,f�\�+JT$�̑h�J�ggj�}>%��D��CSJf�>�q���3�4��};$���8;��F��˨-i@�^L/�{��B�Y���Q��*������zj2$؎�#�C����l�4�7�0��ǿ��`�h���-J
L�.���{����t(��/V|f��T����ִ�$�!b�vJ���	�a�4k���0�О;C������@�~�5_HU� �C�+ DU>i8�I��!��;�q�'�xvR������[�:ؑ�v�̬J{<nY�7��ޯq\�L\��f��1[��
f��5j:����\��B��'a��v�J,I�g�P��oR+��?MC_z�g�:��zo[��]P��~f����(��d�Ze�������Ypn��v[�mDr|�'
�a����~�bUk��-���q��R���p��9҅Q���h�H�Mqը��|t� ?ݒ_��$�&�
8v��P����R�HL�u ��;��G��as�v�z�f&B<ﬢo��l5F��Ft����L�(�<���V�J�� ]�>��,�<~K�tSt6�7�ҡ��؝�K��A ���������<v�����L ����p)�)<����=>Ţ�$l��c�|���+���Wqmf}�H-����%}=��e���>��UZ%w��"�>SC�8�G�ZcD�����#YS��~�"y�(P����.G�|��vA������絼>��0]_qv�x���QS��M�1��f�Ӭ�p\���Ey��H[��B���|���ݷ������T�W+�v*�,����]��sr:e�9�#�Fi�Mq�V�#0��1u�\��sC������9�<!�߫��t^w�.Qa��OXҲ�p�@?��R���6��A�W}3'I�'��J�F����ݥ�[�ȉ��*s�eWh�k�txMZ���gQ�x�7!֟k�u�e��ZM�9)H��½��p�l؟���o����:�����zS�A�эg�I�I�Wr=n���ϫe\�N��� |�_yuD�@!��?�����%
�o[��m]@�~���RK�#���R_Ƚ	�im��׳_0߄zE�\�����R8���O���wOË�A�W�`�_��%.(����7������m��< �w'�z����砡��f癝S�V*l�gH���0�^N"�E|����S�9B��UB��n@�
˾v��,''�%�,��nbo��rz���v� QV"(���LՀ+�����/
�jv���Fq���;�L�=ŋ,NG~��@i�3>7�{�16���A�t���=�W�^���z�l� ��^�����I�R>#�Bz���R{ �#�M���1�+��;�-aC�ҳ��������}`����|��Wc����(A+���l��*(�J"�qN��q�؂�ۥ������$e?;�#˭�ƥ~��Z�����^b	�x$Ҋ�'e:�2[��x��%qt�����*fT��g,{xn�P6�4d_�5rVW��/ƀI��*�y>� 4�?��G����b�x,gO�	�7������T�����l���d��Ñ�W�2�C�Tf�5�c�#����;��T�E7k*��fҝ˻E�0�+�I�q������9�&�X�J�s0�� �ʙv���� �c��Ou����7�k|x��uJ��_��!Uǐ�㜈�(l�|�HN�XE ��P᷼�e<ޑ%KJ���(ƞ)����'�H�4��u�_�]���:ql�siޔ��Z�i�w����W%�E(@�,�#��uUי�;9��n�6�|;�y�
��͙�U��:���_^�=w~���4�-���_s\du�ٯM.�#��Q�l�Z''��-Q'��M����%L;���<Y���Z�R���%��f�T ��4KC��mK�B��� T�&OmTE�R6ŗ���dz}Q��-��H��ߟ��/���(	�hH���Hh����Sѥ�U�5oΞ5���J�-�t�&uD׺�E���X�l9��j�ˡ�Q-��dc��7����4��k�� ���F��QbZ�?'�����{_�n����:h9��ш�H2<M_���A1&0R𰱝I�VCP'7���'"z�@w���O��X"�	������:�	]HB)�K�;s~�Ł���P��Pn��u�a,�����x����+y���o�ndP:�������d���l�>����$���4��3����bi�^K��*�a�|˂��2���U�u7LnK+V����l���kB��S�M����(Ԏ��V��!��|N��;~u�o�!M��x��g �]�n �!��'G��R(EvJk\��	�c�q!Y��9���
G�ʗ��d,���MM~�Lt��j�Zp	�J�z:�@�� c�F�PW5R��6��"4�����_z�}Vm0I�Z�t4�EP��B���7���Li� ejϗ�!�Bd(�|�0&�!�0K��y��#f���'�y��I�/E(�6����+�G[�����D�VBne��O���c�,��M{�OhZ�u
Flw��Wj �+	E7��`6�u��Ip4o�^�c}��c�4R'����Q��T�U8^��vat�'9�0�c�o�k��
�'������e�9�����L�Ì�^�f�(��lp2����������x���D��<��.��m��OLiAd4�oC�~����
��/�糩,�_m�نr�Q�IZop, S9�a�]�ٓnI�"8�L�<v��c��Uڕ�cU&�Ma≓S�όQ���%˘�9ޱ!�񅧱�_�bd;�nzK�ޣ����/�ʎ��0����j�2�y~-��_� Iҟ�z���
1�IE��������^;y�B!@]��߼� {8a���ֻO��x�x4p�`f�3�`�[;��&ت��D�r���zf� ��E����I������YӲ���5~�D�L��ѷA�w��Bx���>�(~B�m�>Z��ÇW�9Y݋����;�$Xo��G����Ɔ��h#��vg(zAm<$��id�lI�5$�ˣ(�{�*�wQ�o� T�{�zsT�;��O��^��w�zOeU�b����p҃�����A����L2�c/�Rz�ۗ� <�G D���`��A�B.�_�A�	���]z��&!ۣ׀)��<VS�������6�Ž�U�g?X
�줤��;ݔ�>(9~��-���Y��;�~��zQ����p�m`�Q��>�:�5AٗS�>?�f�-��A`���׸���a��#�M=�ŉg2e֪��r�Xa�J�	x��_vU���3;=�3�M�oP��|��7�_@��U�E��Ԧ����6�P�!�F%��1f�X�la�-��V��^��)�����};S#����h�����U2�t�P埖MY]r+������Q*���X�>��?\�bq�ۆ��Z�^꠶�u
<iW�T{$,�9�lԳ~ք�7-��h���<���_�jеf���z"�D�8�}��U��<�}`���7��0+���:��0�͑ю����P�L_X���:�#}XW�*.���'d�a#2��שǵ���n`��c"R�L	�U��L=1�X������1|g9�i�?w�W5w��n?�<�0	��^6�ͫ��!؜M�H����s�:��.l�i���SVp��$�r�[2�c�������)����J1m��ݚ4���BV��ò�
�g�'���ע�D�W�z�h#��<�\��)E�r�J&�0�z�::�ZU��?�Jb�p~��:ݖ���-%�<��� �� �={�8���)��Ǣkv ۽���ӆw�����%��{⛨�]�a"\EP$���&
m��o����F�}���4TrW��Gu1��j���p�"-]m��	�s���eP�1����[q���-0_P�Ti��}����>B��Ԏ��Ѡlw%�0�i�ߙ�:)U��K��`��ip�I�P����,%�T�x�ې�(�#�=�7�H:�TQ�IV�7�v�E^�u��y@﵄��9�T����	���3������m ���u�O�?ۛ4�	��_BY�MoPŽ�MǬ��&!7�;-7�r@L)wJ��)�
+F9�:��IvP��/|z�-��v��<�xߪ�A �QB�6���� r��E��3S���(o~&q�m	��J������M5��\�t�![�iTُxs�?a�ώ�?rW7yQ(-����n@���l-�W.Q���|C���7�E���k��k�:j�hp�&!H�Q8�b�Ġ�g/?<ѠMRr��i�����_���Q��U��R�Dp�NN�����nV��S>��p��++"e�X�pv��'R���=?
��qA3�~CR��&�#�g�@��Ѩa����ƙ��5���׽���~�I6^Ϧ�PJ��Z1��2tG]o(}4�_ц�����Yy�T�v
��W��e��t��ܟ��B��G)�D���A2�)�b)��E��}��C�-H����9��
GZ�G�s�ˠ�iם��r&��ݹ�����$��Wu�M�"S\ާ�Nx��[uƆ�ڠ	����F�d������}�w���C�Y��l9+،Ŕr��z�s/��tnΥ��ţ���4X��㵏��fnF��
�=7��'3װ&j�_�H�u
��Z&bOI�����x�u�ز�����Hʱ)bO���+�Hl��$���Ϩ�����?(�([{ւ�ڪV��jyg�~|����V���Q+.�� �SW5���?SJZ�\-#>W���Iv~&g�U���h��|���T����	�L&	�J�>���&�΅vƋ�V�����5�����[�+�}ٰ0o	��P��D�~%��V����s�C��k���r��ͳ�~��/R��L�.
ˈi�ac