��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#�?�l��Z�F3~�Qp|��:��pIۄ�d�
��&��Ađĺ�M�����2�m��ahdH��I�*2L6cB��H��&�a&�sۘJ%�b��T�f�%�Kz�-�����DU���<B\֕W�+f�����o�l�fm���v��W��$�����L�,t_�Ȁ�<�Vz�աW��I��-u�UH�q8/�NT�a;�0��zH��jM�d��}Q2~�ɕ�M=��aF�YM��QΎ�SD�8��fG����V�۵Nu���0��S$Ȃ����XIE�(�Uu��8|�P}"t9̴�ѽ3OBe���Fy��XB&�m��U�!��"J���x�_�+WAXv�i�3)�@��=a�(�H�F�>������E�ɟj�T}e|����%^�F�LB���jׇ9�2K��x�P�v�&�k��RS��d[����wh�U	�7uZ�|W�7�j�PG6X&U3F�б<�pX&��{E���������(�9���r��gv0��y�fk��X��K	B�&i��H���{���d�6#��M���v�H�|ϝ���j4з���gK�՞�3���Xs=6f{��^+�fxnE�o���P��C�# iA����(����m�w�	@ӕ* ��e����[h�V77�'{�0���L}wF���$Q��v�����ٶ�{C�X��[�W��x�n�hZa~fN�����)��9]ؼU/Ia��3ia�v�H�B�90JJ�_QDv���J&�92�uV���\�hoW(���/ ���� 6n�� +�|�{��OP,g][۞�[t�w�t�-	���;�b��5A���<A{��᠆��g;E �55���-�{V6n�gc����R�d�w|i��ૈqK֒m�l�k�����N|r��p�3��k�,;��u q{ L:e�tm��&�u�ߏ�]����z��v�WX�G�9�0��9�-ܩM"ܝV�[�t����B mn��HR�č���5TN-�����G���p�I�p2� ў�5l�m��@���;Z��G:h�30�d��R�Ց��;�)~��ď?�;��1����e/� b���H���k�AfJ�:S�t�$���g�������[
��θ�[H|5�d���fك�TA��� �U�"Ӳ��/l�� <Yp"BN-��~�d�wH�Y(���S�u�1)[�˓Rg�4iuߡ-@��e�--�K"�C��6�㨝}�E25�o(/jr���Ij��;��7#%Bd��e�`�9x�r���O!:%zK�.���O�jV�A���"\�&��H]��i��k���'�G��"�S����ἂ�~�E����
ެݕ_�>��ɔ��!Ap���;�8�Ó�]�Q�I��6�_>l{�	�];��g'�� �C1�g�|���h�TP��F�o�~pLH����n��H�jpY�����sM��L�;�b�}� ��LP_P�2��VP�`����]O�b�e9{<u��W�|�����=�T@��>�;R�;_���R���@������\V�Ծ��8���2��7
�0Z �ᖖ+~�ܘ�-�]�폈t�j_䇕�Zk5T5\���_5邤�A��;��!9!����Up��l0U#�e8Lq��.Z��ܛ#����+�z��6YؓS�B}��Q���4+��1N����Y�5�IS3�/�wйY�A�G�Ӧ��
�1h
���l��5���7OH笚�Oq:Mu~�$m�Tok���[d'qT�aő9�C�����`c �Nb!��a�A�E��V[�vrʡ�����m���9�s៥�����Ca���%��+��E|#q=����@��f�>�z':��}U�91Y(�W�μ��oH=]��j�`��r1Bk���V�o�������]��Ѧ��ܓ�Jl�����Y\ #��	���H�ћ<ix�Q�H~��1lΫ��ݏ-����7i�_\@�H/92ށZ��_ l���P�f�ԋa�nA�l/`��4���q3>͑+�/��#�qKچ{��XF�elG�{�?����=]�1`F}=���O��`У�{��k�7_�g���i�F��GNG#���*
�Zr*ka��Uo۾�X�@`�p�tAsA��g�B�|Ci5����I��C��3���Z7,������G��5�BCr��A�#���1y�Tրf�IUy���hJ- ߴdx��:xzG٬���h�w���f�Q���yL�E�DtY���&�9��V\��	� ��-r��VO0`�5Q	�o�� 7����TD��7�*&M��A��I�G}�#��]�پ.�6��.q�k*����@O)P��u�^�4~YBFF��53���[GScSN�aMy��6��J"�^�[X�㕲$��R��29�P��I����=Kd��&��Oa���}��b��$��=�'x!�n��b�5>��o���@cuW5���T�7q^�%��A[i3Ϙ��ػ�Mw��c�w٭��7��S��ť�7���y�fL|*�?���S�j��ڦ�Dp�Xh	žL9<}�B�(�lFM��C�*M2����~��լ�FG�?H �k9p�mN�	�)��t���� Գ4r2��q�A�-:f~�֒j�I����-����<��ƈ���Y���(X���Z�u��[A'%��J�w��L�6�c/l+փc$�Dq�NdS�a�A3�v���!�����.9�kPX�#�PxnX5��!�;�+�pt��:>���/p��l�nb+��{V�N�cDsY��n��D[8j��n��I`��C�N��XR��?,:��=�ζ>
��/��Q?�4�����\����H(�F���
��SS�]���<%l&l��`;W�5S17�D9�"�hъm��4��m��.��8��+��ƩA���b�Z��Z[R6Hl�Y~��W�ʮ;�t ���`�������6�M9�/ [��l�U
$0U��GA��,T'_�;Nw#AK�(�|�<^����j��i�Y�F����j�I3$mN�=���խ�)8&*�ڂX5*��G�rl�Ҫ�@���S%�!%���aг��d��kU L*�{9\4��ሆ�~o�
3�q⾘Z $�3K�c�M�1y�j���X�I$��h	O��-!JH4�t���[ ��?]���	��J������x�~e�I0�9�H9nh�����Z�R���뷺P��l��WG��ˮ#kO���=�r	��g�"{A�Uwݦ��%��ؕ�? M�fyI�X�3N��Q����{;��Z�=�,]"��10j_�
�+���}�F�5'OK�h�2�@Ce�)�q-J�����s��<2���IE��O}Fa�@�!_���'H�$�����zi�ξ���f����F��3F��v�3c)R�+g�DGa'�9ϳ�'���u���C%҂-���~^Ag��c,�ٗx��9<=�ߩ�����>�7b&P�]��\��p��5es��-�]�+(�䟠޵�ZEIޝ�ϸRA�a>\F^B��<h�������9���,�������ǂ:����#ɗ���3�9	�b��d�F�޳�#�զa�ø����� mR��-��]K�0��"q�n���N�R��i@�J�]��`P�E�|>x�Y�g2�I����e|��7�sh����t�,��c�t��ĥ������*xC��04�H٪S�����a��H=z����I0��<��o�o��Cb������ �(@=���g��A�v�q��!޾m	.�V��rH;AY=7f��?f)�:��j����]�=����.Ex ��H"H�����9�&�P�kϯ�����z�ۀ�@�VnصS���a���J�2*TL�����V�YUF �����F9뜯h��3��k�������[րԹ�b+�M]튼k�P��~���@��8��~#L�륮p���E`�ϸ��K�zJ�=�C@�]ͽ>��n#�BX���-P5dL��CxAo���|9c����d���./��[��?۽)r���|�h#���Ah����ٶs׸�q�#U��+�\تz���<B�Eg�	�����h\��7�>�%m�Z0���L\�P���@.Ck�� X�a�!��Yp����2��̹�i�ɍK�f�����7��Ե��J'P�S�a@��PwG��`A	$���%WR���3�{OQ&����'���4ꩯK�J�^���?����b윳&�(����CiX-ށ�rC_6�1���W)Ȝ\׌9���O����l�񝒋�$_�q�Lp�����?ۃ<�a�W'Iŉ!c����z���WP�V)m=���5�7Ba�b�:�B97i����5I��K��VM�v�c/.�v���Tpq!|ҳ��L�`ۖ�7�c�Y��.�?E荪�A�y�I��i���� ���R�px�ə�2�q�e-��c��ep����8��`�.�����ѱh̖�y�V��X-��et�a��WB���΃iєy)�]��$�'��������E� �*�t�N�,!}�Q� +P͛&�+/�v�K֜:���Þ�#���&�q�4��ɩ�Rf�p>��d(�a�p����-v��z�R���@��;�)�����a���[�sՋ��h��h��*\wǧ^�" �}�ڕ�Ӓ�{8���d��0�A@~��0л�\W!#-Q��+q�eع��o�	
����푀 -��Wʹ��$6D�&�F���������L�cS'�9�XI1��Uf0)^a!l ;���1�&�μ]K�Vɥ�|o�K�ʖ����S�ɚqL|��E!n�(t�!����p�ʾ���ƴi���t�C�A� D%_�E�63���64�XDM+5e�\F������O���!����lY���ԔS�
3��@G���B�CQT�AdRN$'���-?뭯h�}�#������b�ե�h}��ɝc<�yH��#^Fu�f�"I��|ֈ$��4��/D_�P��-����.���w����H#��Um�h�N1+�H�z
��X�m�r��:r�R_[`S���\�V%F�^�_'nf�TI8�d!}��9�ĩM.��&Z���G�1Hy��ښh_���_mI�V�%`7���>M"����ռ2�i^[ͬ��h�¯0�� ��6q���V��}v9��-�ZOG���ӷ�������e�����3"�o����So�Ah�q�c\v�N;�:4u�o�4M�0�@��l��N:6a�/��E��o�9�d���/G�W�c�0i>���n��eb���.�����[3z[����7��9dX�,�?8{Ɇ���K&];�>����L��L',�tER������	j���s�Ϯ��ͬ 2uO���[�0�E`<l�@�H2�m����d�{*E���u����w �P~eI�Ӎ�B�j6+�z����8?tPe&\Q�5��!�~7����Sv�|D���-�!�<�8��4�	&h|�d�Ŷ�^ɱmD�'�YҚ��Sqh�i�'��CVB��4�A�SЂ��ᑭ��o��e.,�22?yރ��k�0���6ڏ��Я�������S�A� %;C��|�W|>�2�$t��E��dIn�>[{=py`���q?�a����x4�rnX}p��pÍ���z�A���W�h��l�J��O+F����y����b|c1W�e���C
�GFM���� �5q�ʂ��B0w�j�����l/��N�&I�F�<��o2�ɜJ�;�.�u������U��l��HE徦:NA�f�����Y��R���$?�>z���YD8:��k{ۧ��E=�N�dOs˵��Ғ��$�fI4��sZ-ӽ\v���*U���9�z �ubD�����^�C0�0$�%�̒7r�<i�&�F����¦��jC���2fĢ�q�]��\hJ�÷b�	�6��&>�.})Do^b����l�7���Yq�)-���5"���[-6�:���,@*���V9��Ex�Q7{Z�2���B<M�z��iv�7pXU� &-]�%Bu��@��D�IB��blDK�(�5H
e���Р��T O*�����`�'S�Ew�VC?���o���<��+�����еZ�r���C����݅�rݪezMs��"��hÚ��E���IN�`@L�锩���bÚ��.�̧7�OI&2$�>#]��2R3P7��MU&q6 a~�]��X��J@m����J��ln�ȵ��n�K�8����<jF�)Σ�W�,!��HQ���]���wY�$
j�H���P�cI�;g��]�F��e�su��%ڑ赨	�F)Sq�Q�P�w�D t�:�!M�
�'M���x�-���-5v�ņY�f&V5���}�Q�$�s%f �f��&�����Ghs^Z5Wq�/O�5qa���yu�E�p�4��Js_:$��3�N��F� &�:�и�@��6�a�;�^Jԋ_n!c�*����#m�E�w@q;Œ˫H�����H�O�g�ӛy_%��T_Jq~�Br躧������(�|�����b����r�)%Q:�9}밞Mh_���j��uv!�.��D����������ɿn?�>�nn2�Ns�4��X�w&��ث��-cC����h��	����X*)Ԭ�.*�"�>��Hq޿��>� ( ѫ=��������%ɣ|;���	��$�;.��0��b-�a��?"���V���,�cD����o���%�H$�v3(��!���B3�� ��biS�~���w�y���X:BA��"X�^$�*26�d>J8��xg�p��"Ã�F0.��޲D���vv�A����o�n���(/W���0�]\� gʣU=�Y�����&Kw�.lk��c؉$���+�]<Z�.��"���*H��b��0-=7I?c�:H���'ڊ@��5X�5�d1��1k���%���3��W��[q�:C92	��S�����b{�r�� �u��0/G��'�*��B�V���7���c���� �u�O!��bcR�x��Ӡ�zx6 R�P%T��0Мp�?p#fU�;o�*�*��)��1�&�f=9-��4��2��P"�lI��a]�@w;j�򐕍]�cQ\Ŗ�|i�U�@ۂN+A��l����e ��:�K3��$�oM����u�3�ӏ�`5���M˄��R�`��"�QX/�Zĝ�OyL��20�ݒ�ڍ~o�A�+���n�k���Y7_�^����D��m��M��,�G��kp-�
�
j�#��J%
9�mvaI�ǈ��A��7����V�+�f�����e(y�n=e�%U�iҫ��آ�ASel´�4};3Wd��JTK�k�;~'�v)�L�.F��P9N�r��9b��zoW�\�v�nH�C�\Eh Ɣ��ӳ�CT��k7~o�#����`�Ły���5�v%N�tCi�}r6o�@�-�^�~�2�(��u��7]���i�h����	�9<�u�GA��1���
��l�O����-d������]����+%�0�V&z�t=伕�U��F�Q%K�D��E�U�V��聯��O�_{ww���)T���c+w`y�R���q�Nw�;̌����tv|<�3��FW�.�5<��B�gm|�4��C�G�@�$6!�(i<�c�d��nt\���������?k��]2#�=F��&��������Q�j(5C*t�bʹ��?�-(��xQ���W�,�KX��Kҁ�_B���#���|�x?u��!0ʧ�&*�m�7Hy��my�-$C-}��D���<]�A�/���Q�9n�B��s��_��!�+.Y�2�e��V�o��`Z~=���	�Y�H5�ND�*�[��q����s
�Rޑ� �	=b羔����U{7y��(PL�����8AZg9�S�#��H3�����Ķp�I�]�3�3c0��k��k�
�ܥRZ��	�C�#M"���CuG<�=wAxF����cG�'�~ɥʙ�Z��uk?��⿨�1��ɌL�;r�l��y0/�����=<Tt����6���j~#�d��&B
U���g�ֺ�=���),h�g�L��}�n��/!��N��#vTG�('�{�8�C~MWv�A���(��SEaa5�'�M����k�ؠ���ԉPя�s$ՙŷ�у����7!��S;Z{��0D$���2����S����D~c��-.T�yIF,�[o�ODu�iO.X<ȩFA�j:6��O�&�|;{�w��Mm�Q}#M�V���:���)�uB��I�ut�ӎ
��0w_���֎�!�$��_�'P�xz�==�_y��Yd���b;"d�.��Ǟk��x��ڟ���t�ᵅ��*��V��S�4����'�\�a8V�&w��[���������b��ဉ�3���@��'�=�<�:e�ku��jZ�C��hN�D-]w"�#s�h�Y�0<��A������d�֮�Ǆ�3E,^ #d�d;_�U�Y(�|��#f�ǽܨdG��F`'��t̖����"�'8�B#њ�Z`����+�>��ѡ=~�w`B�"|&�g��F?%K!󫿆�7���w:�6�`� ��W�̓cr��c	3\(>eX��:㋎����eBɽ��4a�a�,�S�Z�S��V�#o����Mev��ь�_r�pQ1�|u�Կk�a�c��u��8�}(�kZ������r���`�f�m!�i����rZl�y&yj����P:d>!Iw@͛��Xv�S��-��f��'7Q�$Iu�#I]�nVΥP���;��7LRi]��.S�d��ԅF�BWM����*o2�yۜ�'Nԇ*��zx؜۸fȨ�Q�#x�ʡ	����C��Nq�㭸E�'5��&ח���n���.�0�[��:�o?��a[V�0ф{0Z^SOjl�,^�+*���w��	�K�J���1)Z|Ƚ��](�Y(z0�j��Q@�@x�׻ ����W��87=c ����3#�<��%G�+1|�hvm�\=Q��1��o�z_Z�IB���~/���n	gd\�Lq�q��14'�PkѼ�	����Pq[nx���g� ��Q�y��-�l%7'��H��{�6��p	$���e���S�}hΌ�*�T2�2'�j��5�����T��� �l�(����'�:��X/7�8����V�2�:�9MgŧF8���kz�O �0v�0;��>A�д�0�}��,{�Z?���x�cLx�+�I)%%�u$�ț1��4}u�qd��0O��2y@ma�t}W(��/88�����
��2���h�~ \�\��j ��	��U��޳�x�Jʿ�w�$De�s���#��ݝF�)M�v^66�7uٹ��r�"X�J��C�`0�91v����!���fu�|8�&�/8X��s�'��:�y)��qV���v�l�;�Q�x��3�ֱ--x%z������G
�+5���k�_�X��y��<��3�C+��h�d���/~ޞy�-Б�Ǩ�1}U�>è#SBis �l��i�M�r�z�v�_|5-�dɆ}f�����W��M����օ8M�7�����O[�^"s�4m޴|j�%�ʋ��q��pR?��n/�1O^�C�<�;Z?D��rz2Ⱦ+MT���lM.S�/݄�/U��M!t(QQ�p�kv�ǝp��Σ�������$�}�&N�8u҉L뛼\<-���;/��9B�����t�8�P
�tH��c�r��u���/{�@����]�Ѥ��!X�����siֶ�XY��=��g(*���[���I�xO���J���2��d�Na�8vVh�QK�8Rh��R��
�J��t�m�Si�hw�3)�� l��\u_Ҩ��<�%��+'�B����C�,J��~C��Ǜ5Y�m<�O�0�|K���|� �pSQ�k˚���'��wl��>������k<�s���P��E��K%Ɲ"@�@-n�%�}E���%N�ӿ!�c�{0l�+[mA[�5��S����������Y7���b�|�����Ȇ)^Հ��P�K����:��B�me��F}���ڵ�3��=�S����d3X�2D�~;W�W�'}����ZU�ڢ�c7Y�vU�\o�w�P*��ǡT�+M;b�`�=�ۃ��{Ls�Px�����S��ij������ao�B�+�]�oO���mZ��n�x�M�t>�AI�%h)�_�
i���2����O���M)_��:�2�('�;6ħ�
_.�3�,z�?!E"!d>J��d@��H	�c�Үվ����es�H�Dk�7�lT�ϱ��!�8���f9l��v���6�GEA�k��G���,�������<�-�+�ڋ����<�ְE{�S�:#���
���.[��P��e5΢��^�{��]��į����b(����K�u;}��g�.>/�v�W-4��8Ȋd�p��d��;9���(�_Ϙ�dWpi�2���"{ᜬ�bY���j����"��,���:m`Ó���B��Ӄ'.7e���%"�Ը~M7�����.����@�Ea��=Mt)5�Mauw�˴�����L	?��m��i�/��ZF�5P��T��d`�y�G�0L\�U�gX:t�0�Iw=��uc���T�K�a]Nv�Q��d��:
^!(�>��Uu�H(��+ks��c���%e./�#o�2:XN���o_�(��>�vRt��q	�����ְ:5G};����~���`P+�uOKJ������S��(	<o���z��~A��g?��-�"v�!�`�wu/�݌���4�qi h4�ao��S1�G�>t�:H���P���n1>��T[=p���Ɠ��
18��c���b�����-o�,�5����_7 j܂�|�! ��n�1�Ub>��oƛ��)�ƓZ/��[�{����Aw˙�I�}�#ƀ� _���e֐w�OR��D}�B~_��Q2ԭ�������>(��ϭ_��������S�4�:�C�K�5��� �}G}I Mk#����Sa׺��r)ݚ��_��1���[�p��L�-M�>�����I���F�䘋��'��ᵤ��7�i�w�q��޹ЌxTWY��