module compress_tb ();
reg [511:0] in;
reg CLK;
wire [1535:0] out;


binaryToStr dut(in, CLK, out);


initial forever begin
	   CLK = 0; 
		#10
		CLK = 1;
		#10;
end 

initial begin


$display("Starting LZ Compressor testbench test...");

in <= 512'b01001000011001010110110001101100011011110010000001101101011110010010000001101110011000010110110101100101001000000110100101110011001000000100110001100101011000010110100000100000011000010110111001100100001000000100100100100000011000010110110100100000011101000111001001100001011011100111001101101101011010010111010001110100011010010110111001100111001000000110000100100000011011010110010101110011011100110110000101100111011001010010000001110100011011110010000001111001011011110111010100100001001000000011101000101001;
#50;
end


endmodule
