��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#�?�l��Z�F3~�Qp|��:��pIۄ�d�
��&��Ađ�gڌqyI�3�F���i9�G���S,&�׸#����o����<���?�O�_3q>UM�|�����}�}��oE�艓��y��%���t.d��Q��V�yW�]��gә�-d~ͬ�!��T�-~����5�[�����Ӌ�:�S��"WE�|h˗ж���c����<���n�xyc�O�%�j8Y��.�Y���U�A:!� }S��d~L���/x�ؼ�['*Z�oɶS$4��h��iy#`F<Y�Ft��Xu���g&v/��Vj�%��3 nK7ȏ�G-��H�*Yƾ`l�fes�{M�9�F��?f�+��p�"5����L<�k`�o@�d"?�KL�G��N���/xl�W<�k]I�XJs��+	��ĴJL��i�����H$y���=�ԙ8==m����7��kS�l�P����,���
E��=,���:f�)�拯xH�ٖ����J�_���a��㛴n� ��xV7���;gY�����!���
,��k�w��Å`Y���{A�;E�U/k���Zc$*����������A�[�������Lm+�Wu�Mڔ��@�9��F�v��@Ä"ܖ���e��Jr��]C�8oN�K���-\q�PuEJ�')��z�J��A�dѫ��cw�y�O���Nrj#A�n櫕�ۚ��P|�5����M�6�y��ڑ"_��t@�ș��{[��E?p���u�ֺᵃ��(��ؚ
��kkŢ*�g��:'���	z�F����.�s��\&`�E����!��;�#���v�����;��H��\_�]���5��KV��᳟�^�@&j�.<p�e)�f�7���ҏLϧ<^뷈�>� �J�8R~4H��N������_��L��b��	���b�75���#�d1Aί��E~��L��X�Hk��Q5�j��r"����զ����T��z=Եw��t�|T�K��Oq�Z�E~���}ʬ�m�����Վc��,@�yD���S�_)-;��/��ch���w���EJV�b4��щ�!C�'����P���Pk�dI5����(F��Ž�iϚʇj�q�����7d�!�T��d�� Ԗ�6h�^�)�-:d�4%Z/^���7�x%2��[=��uk��G�7���2��������5�Ρ٪=J�![N���s��D��F��F�i*����SJ��b3y����8�5��I��lN�5��n8�I�9_A)�?f��v��7-2����7{3r�*̇S W�%B��A<	f�uA�e�>r�xza�K+fV��9��8������͟� ��KO��"Ԍod�0vz�8�4t�o�	���|�Y@tx�����G��Lv��o/�6��v���b\�Ko�,����s�g	��t<��۵IZ�B�t�X{���ΠNz����m�(��9*t��o(�)�A���ɂ����0K�j�hz�r����V��k��?�jY(F�P�cZ}�w�be!�Y;%�V�!1ss�TR�Gd�m"x�Cy5�/snP 8J��2�/H���'�7Z�͜��_h,����X�i4����j�L����ъ��:j|����#��mo_��Ӆ�� �^�"��(?�A��k W�����\�ZH�DK�|Hp5I�� ��['�N��7xU�d��#�n���S�;��>�[y��`eX�d1"�I62AY�1_�ĊZ��A@��@�Xɺ37F�H