��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`��T��D*Fd?-��+.6���L��[����4LZz���aZ@�Tt@��8���ű��sY?��>��
���351�|a�v�"& �o,���!��cze��y@/��#�	�M��-�I���C����a���
�^5R/CrLݶMqL�7�J�)�e�N��
�`�u�u߳��4{� ��Mrƨ���0�,lG�����O��X$'�/�jɭ��/�KfxF0
brIr��V��uW�.�z�vτ!���Rz걖���)�Ӯ����^���X6�E9?{%\h���x�~E<�L�=�"&c�w��9�[���.I0��A�Z9����$.�#��~�Q����ȚN�����9�Ö-q'�=�����%yD �,�,/����l��r1�ji���d�*K6��=����� I�v�HڞY�Q6�����U�Z�ֹ���ʠ���"��$d�p�{�۝���4x�RmC���wuݷ��\�]��Vh5t�����1;b�~!:���a,zi����:�{���|4����v�k%�f���G��E^P���}el��]��S�����j+�Y�'(�'R��@ѡ���M��p�UV
OnN9r��|�׺�X�F��{�L�= 9�ȫ�1��0�(CB���H�M��`=8��u�����x��^�XL�=xM/&?�����HR�ϩ.l/oɓC8��zé�ySD�IQ��:\�S�Ab���Q�����9���X���J�jnW��~�8�s�$A�J��
���𴒎m,Ue�.���ym6��b3�}[��'�z��B�����0Ђ�_��B��ﮤO aˋ_[{�Ѝ	l������&�������S�%�l!�Ϟ��7S5
�I^�]�3�������2	#�.G�ϴ�Tvq��h;o��rd��S
���7�I��F�'D[��?�y|��Ҕ�����
�T�o�7:B+�Y"�ڍ����N��J���A����3w{4�'^�4H�~�$���ͱ��M30y6Iݾnw���/���<Y(ב����%��R�%�����%�{1ז�7&�����1���,�X��Z6Ji��{vQ���q��wXЌ'G�� �����J�0ض�HK|3�O�i{��� }���xpLr0q�Ѱ�bT�b2NsÂ��9�%I���7c�=p�ǧ7�����g-�s�~���@�\�5I���4�����f@[5��1�dg�eaF�Ց��W}M�L�6�vը�C�G0ք�����%����Lw�)9AS�kĽ�i��_M��Y�$�#���uȃ2]ߑz�pJ0R��>:y�qN��v�\1A�=˕�hT�]g � ��|�PÇi���Z!��n���i/�Jj�.��Y�!�F�D��� +Q��X3U��ثp�@�	��C�_$�+�HQj�[멋���Sw�	��%'�!�ȍ�P�K�FzU��B\G	H�C3��ڒ2�h�\���<s�V})-@ۏ?gO�'�Xk�_�T�$ųɋ�R��o�x'�u���t����㓢�R-b�����	h{8u���9��+#1s����7E��J��ՠ*
{�V{�΄,U�~�Ve� bf���;b�V�B�1f��G�}��z�}N�F��h%�a�g�%�*$ą�mI��2��,0)8�54��?�����Vm?$�Y�w���Q쳰�`W%�uEHi��Y�K,mzk������57�D�[J��$H����L���]s�����D��EM<����m��9X\����rU�	�jM�ͬ&4hN�5��;��)�tlV.��n��h��R�u  �I�zt҇���3�릦�9����e��e?i`fac
:$>=�@���F}X����-8Ka;4=�K��.�j��|��tFLP ��Ih\X/��1�w�����+��ұy*MGԗǞt�ˑ8?���ZA`�܄�ʡ՘9��ـ9�D���t�]�������u<��P���2/<��p��D��'�"���� ��G1����J��7�m��;�8z������X�qt�?��e�[���߽��D�E����'���O�.s� �;��?�<qn��M�/���(��H�E�22h.��*�n����)CW1�����:u6�\�|f��#�U#\v�@�5�q���U��F��J�)�t��k˂>�v�K~�cV��l�n=�Y3�`���+�7�����ʗC���\L��a� ���r~cK��[n��vYK@��^�wq��g� ;Z�H\¼5Gz8���z0K4�,�����pNT�ũ�~���m�J��;�-�^Z���������o�4���f�l��㊲󫄝Oj��'�x��cZ ��3���$�Q�|N�?,y9+�^�Z�u��(�f~$�xvrT�a6QvA@]����#�[� ���{@�is��BD�NQuw��a*��cNzã�[N-��ʫ�$��L��P�O�RS$��t�Ĝs�}���j:��
% o}YN�_���=��J5��}h21K�g����4,6���*?���`��2�D��'>�RY.����e��PJT�"Bv�ŝ�&�8�q'T���95B�{��O8����lL,!�j b��rˮc����ŭJ�-��B�_�n�M�j��8X9��l�Fc,�j��ɓ����P��)τK�{�g�7NL�a'66������:����2���P2SBj������+A'kpX�9@A�$W��-�=�oc�����4:GL��v�����?�8��z��T5��/�Zo7� Edj�N��������Ct���7b� O�A�k@�,�6�G�ٳhX0�k,#�sB)���{