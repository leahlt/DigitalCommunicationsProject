��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P�|5js�[`F�q�t�(���(-jp��
�����-V�N?�;�� S���H7L���S�w�Wj�K�DP2�_K�=@�%��՜��-d֥��K��8 �R��к�u̧J�'�U,��O!`k�	vR:]L?�q�`�Oم\�y�ˆ�a燺{6����/���
�C���2�M�z1S=^�J&��7�}J���b��ĥ����g�S����j�/FY��E�ݪ��f3E/��m8������RTWq�u�AmҜNh�=P�l��"������8��mi	Jm�l5�z��&I\Y	�q��H������y")��o��Ә��@� �rL��x]��z���]C9y��j�$-�zғ�NK���
�F�;|�G/p�(�}��z��n҂��U�S��(�sF(L����wE��{�������#�W�Ft�;����{�͹Hl�8jt�domk�%��]-߃�j�a~��KN��Ұ!����[zn��#��b��v��H���,�
 �09�I-:Qwf�0��:e�#��C���%�$A���a�~�oQ�,1�Of��dBT-���^&+��%O2_U ˃d����m8xO�ፆuN�g������M|$vnA=^~=�A0㩬���'���r��$IH�p���~�v���z�d��(xG��Cue��P���,�@��C�yx�dGp�D��jqk�2�<��SR��ED�}#�)�Q��[��K0O�[x�����k�[��nP[�(��N�x[����C��	K_�4X�Gԍ����:
��F�y�*4K*�J,�9���C�c;��y�*p�䎹i��u����c)N*:HW2*g���j�<0����R=���qC�4Eʊ�*䕿"��m��i���8�:��!�&� Oja��>��o��)gT���.dG��ʬ3O
��4
��5NP�S�&����j��m���%��>�2�n�C�ʹOA	���me��W\z����^FY+ݪkp��1��qH'	�� ӵ�|ݮmCN�c�5��_��3���iU�*�KO�6T��\!��¼�<��p���y���������(o�=��֪�T`�
dph������U���y|�n����J�$ZR �M�Z������L��������E32�wB|��}�
�'�*j?�Hs�8ΜZL��� thCdT��ۅ��u�	(�ck[��ʞ<�F>hK��{�9S�ɸ�1�di�i	�£���-A&�+U��S�H�����B�J�2?�:cqԆ��V����[��g���A�Qk�`g+�w}ɕ�f`ر\�Z�^o1]4����%��ZK�+�־(����>H)=�=���$	ie�z9�[t�H���� !(w�jm5v�IMY85�o���#���bX����5m�"/�v
�ez����<������i:����B|"�T��CWΖ[�
�j��φ��W�ق��0��2; �X�&0YAbA�>x��^G�!.�@�L�^ �b���(_F+�C�Q���b��b�r2v�S���#T�)w��t����m�+
����Vϟ��?n���[�aƝ��RP����7>���d�ִ�8�e��E�&�Y��Ij�y���f%��bIvN��)�|�#e��nC� �!�ZU;��P�ɿ8�V�k�h�fe�'J�˪�SQWuQ�)�%��1hAO��c�n+��rY\�D����bfpH�(?I�o�?(�޵V�d�<�T����v7��7MWx^r���a��H��c�
�)��(�u~�����$���=���"ws���X����o�@6��H��%��H-V�%v��_T�D�'j�b� t����3��]!�,�*�A� ��(�g9p2����{����1�y�f���Z[�)7��������!=��6�2	k��&w�v{�V�|t�B��ޠ#���|(�F}������f��m�}�ڊ
%I˄���+8���j�xJX��©t��j�s�U�4�@nK�4�id���d@���F� 	,�QI�\�.UU�]oC��k�X�i8� ����G��̴B؂�_����k���t��|^�����ZP>�t#*�S�T�W�	#"**��U7P�E���?wH~� ��(>M���={ȹZQ�K~o�D�q,�
��������H�ф�Lj��W:���T�:�w�����&�������p��oR���H���٥�ï���|-�qnIl���v<]uJ����[r�4QA|�2H�wJ�O�G�[���ea�E?�Sޯ�j֎��H'�(�NF=t���v��9��r���ԯ��ߔ;��o"�O�`�q�e@)�o��b�A��N{-��j�_��"6�}�R�`���t4��ݯN �� �]�Cj��Xu�77�I�T�80]��`��Hl�VK�|,���7��D*�%[�O�It���H�[��ӻъFE���Pf�
��ny��kՄ%=;]���8rJ�3'<���65��68�����g-D����N��RjN	3/�Y�
&֙����7�S,��y��{]�r>�hR������7��f���W�I�s�T(�L�o�4�B&6/ct0 K���d���B6�j�@�_�8�R�����u��{����txx�Y
ny���D�Ѧ�־n�����_��;�{�PL',Ly�����Y�-g��p��Zj8�t���LPB�1d����Q�N�7��&2�������t�^*6]B��͛r��h8g��'"�):���7��N�̓�:���:��j�� ����3X"��q?t�x��)D��J�W,&a(G�o�C��3�;��c�ן�{ �ti:��Rrm��nl%p�s�*�v���gHIg�@�y΅�2� *h�J^1;�?��;X�rwm�gf�К���>.����{ �ǲ�1���?Y(�H�L?HՄ�jP�!�jb����e���z"x2����ZJ����x<���.צç�U����O���9��`�Ā�rH�q�-���ث�0 1�`.O��yL��6[M����(��	#�Af�L���0CԔ�#Ň���,(urI��t�o��9�n�g��H�>�� �7��^�����'|�%,rݾnNx���g(�|­{����!��0v��S�M�j�~�a���g��{a�U�P��x�I�$(���Ր4K�O(6�@���6E��3�F��b�P�)�u%��ՌN�td;��,���n$Vn2d�1��I�B�G,�&?��$�5�ύ8$P�����!W
j�H��ki��mc��#��e/rHp��,�� ���޺��q#�y�Cb�٥�ˠtOf��z�Q{p��Q<0�S��S����&��Q�l������Z̆�w���a�:�y!���ѧ�I������Ն+'�4Pf7�:��E݆�´��=^��J�j��WcB������5�E���<-���k,Ea�6@=��J��Cu	"=k3&�'�׌"ͮ#+�x�i`-4���*Qc��C^�6��t|(j��d�*����+}e�/l�E)�vG�;$��4W����=�p�Ib����D�U�L�c_:�<v)w�S��Εq��������Nb4�9��翨��%_O��Ф�����i�[!���`X���Gi��n	���D���ad���T �֥�� ����hfm�с����1��	��e�v�3{�	��on��7O&��W�~�~B`'<���te���-�������6EJ��_�E��'��A�[#
s�~�i�Eʖ �}�9B�(��qm���|���5{Aw�TėG��|U�5��)��Yf�5X�Q�뇛���Og����=�!���m�v��q� D�oxˑ�����N��n�r��2;�S�U�'��>$���U*~o�u⸽�t��!K�G���/�$NxPN�VJ!|�����`'�Ֆ�8��8�ޜ��q�M�Ie:,鹌E墠����	�/[f$;\$R�#��͝SI|<oձ����̳�Zծ�{5
jZw©�guO�^L�x��8�/�u����]��F�ޗ�V�N-hs��q�f��CP�~4�
�
�V8�zl�k�[�z��5{0�<_�b�����Jf���j�'�3�ݜ��̍�������fĕ
2�=�(��+f�U�c����S�o��q����Ld��NC�z���gr����AG��ZZ�}g�����S�� %4�4�$�R��N#B=&��VCb��-�wl��C���c^��C�0���>պaɆ��-��|R��h`�J.%�.�J�Nd��&��S��e�F�W;��U^*v�s�je��<���m�]U�c{:�knA�Ӯp!�A���h�ѡ�P!�D�T�D�,�Z-c�k�2�Vd���O�}.���6op'\�@�.����B"�+�� i�{�չ�+��������m���KpW�^�e�N�2`�+�6]j�{����З�����q��bi�ॆ��s	�蒣1���e2��������m��W�˸�/�w)(�+O�\��Wq���{^:~�y����7�l�R�Xy{<�9~!B���rC'W�}��e���62�kܛ�t�0(�0���Y_לv��{R�<�u��9l����g�o��G���\��l9K7ms��J�(wp0��n,�]�^pܛs������j"���B$yw��sb%켈�Rp Z@�c5��UM�LVA��\�}}�R��|6�() ��^���ǆO���J�'d�Bis:�4p�/Rx�fZ0k�Ib�C�pE"W^�����轩���BU�[8@&�@+^��0O�׼�Ɗ��A}o�5�۳Cߺ���d�+��M���gQ�o={w�{�����hȾg��P?Ф��h.�L��6�ks/#B�k ��?K��f��]�m1�v翀>�B�?=���J��]"��a.~7���Tm�^W��|K�g��z���Y܈�6�3z��P��]�v��"���͉�D��*T*z�AG
4vcn<<>��:E_yV�O�ᜤl��"j;6Z(����eD8u�ũ�F_B��V��Ui|%b0Fn�o8����=�{��o��PE���@g�H��LTm���,��+S��x1]bȦc�m\?���<��6���Rםq<2�2_�jkN^��A�����o	�Y�p��(���݉�N��̑_P=|>X{mq�u�"�����֗ü�C��=I���w85}˵g�Du�k��?�>ʈ��.�6�o �y�e�+~b�킝�u<�;�iRNX�4xq�pf;�g�`�P�����?d�����C�������LS��>Ȥ�N�"�+��aw?3a�sV��G�gE�s�����@�&�<���n�z9t���Owd�⟈!���O�6����l����ٞ붪��r:��j��B�#���)�����a�w��j�,*�^�"
�T �[7�����6b��w(��X:�²���:_�j(�X� ٳ�R#V�T5��J�T���}��[�ywk�{bF�}b���7SgneF������k>��� �&��N���A9���Q�3���3�3d��e�^�e
����yܗ�:0���w���``�z�h��r�K�ϑq�ng_����֘��@#0�Ho{�X�l-��	�mb�jX���aò�v��t��+�@È�񳝯��*������=<co��&�41�@=���l}�v��J�������f�"Ì���E#�IH��<�-��*?��kݸĝ&�D�L����|�[��M��@I)����z�!��yܻg�2q���x"�@�
ӥ�-f=�N\�K�v	��M�S2f��nM�f"]��rjY�3Am�4Q<��vK�n®��]�D�����6���s�(I
�n%�S<J��1��ʊd��h�[Q�������7��h8ЃGk,
a���R�P��s�x������Eՙvڋ�}$#e�$}��i�rd�P뽊;&ME�^ʻ�\�Sj��H���ν �'l�|@�=w�co��֯�LXU/�����p��ݏ(r�L5&��)x|}��;K�Yzb�;\��K��䂐�s��C�;B����
%`�9v}�< ��ն� ;�Ob.��u��дױ�i6]$I�r[!k�cH2����D�s�i���xz��ؔAF����ɪ��4�&�P8�\aZ5�����ΎJ2�U���ۺ�
jQ������Ԩ^�̇{'f?���i=�yf_�����K�R�h����=��u��HJ4��c~�8��r'��-2*:l
!ߋ�i{�%�¢PM�vg��nQ�f��2VD"CU��2�X��t�KY:��l��*��Y�4������6F�hth�ba❔�oE�Ƚ.�� �J�HU��Cx�7(S�U�E!�Y���@����r��U��v3��\�-FMڀ��s�����oԄ.��&�>���Ĵ�ʘ�(�d��1)��J�$�K�h� �l�������(JH��W�S��=$ie#د��P��I�H�F���>��B~�J-�c��><����D�N����`��=�LV�?��FAͫGH٦�Dk�t�\����\�=Vf�w[�Mo�Ɲ(ʚ�H3�mvĎ��~��>��FG�l�Uh��D*�ǧbaM]��:$s!:���W� �t�f���F�tL�3A��.u���R�Ѩ�����&�D�Wix�#�\� F�6}�0v�YUN�&l侢�GbQ�N�	�� 9�}"��f��n���S)N;!{]?��P;��E��@\ɉ�gZ���.0Y�����bb̌O2O����`�`$iJ\��
T"�����WE�3
�2d��\�x<�ז�=�l���	��R1���ƚj"�� �9