��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P����z��{}H���_Q�hФ���]xy�0�|s��9߼L���حe=�3�����Uh=8G%�t���n�4��D�cm��zۜq�a��?w}HC�#u¨�`�L�Cަg
WS�1f�k��Z�WЁ��ehg�+ݖ��F�	Y���җ��2)W��Á$��%��-�B���C|;\�z�8����P�����`��:���\���c��E�14�QC4��l���&�d�2]JQOmFåX
Ѱ��*��~����kp�˴��׀Z_ҥ^�(��
��ve���g�;�RR�Ν��u�!!M��Y4X{Vp���j�o���o�Nr/D%1B�/�[��|��t��w�-�DＴb{
ך�snv���Tx�7`�l�9�~�˺ď?�|��I��;�E�pJ�S��ٻ�eGeWV�[��؟;�ڂ��2���K�����$gG*D^sY�9آ��G�{�-q�^K������M3T��G��PM�Z=ŗ��̱*�(a!�m�6�u���� �c�b��ʼ�:t��� �?�ȇx�&����䗶-������R�5=[-+z����e�B�S� �I06,C��B���Y�����)FPh3e7�Sgn ;Q_K�v�[��+��WL�F1\�D����+Ǭ���}{z�iT��D�k���23���Rf��H������`�0�R����(��K�PƢl����VM�=��RN���G����O����k ��p�^���cL=TAHYړ�J/���5�m�����ԯ�m��n��QX�9�t��<�W����.p��"��eԎ�
�<�Ɗϊ����xk�tź���Ҵz����ťaY9{O.�vZk�d9��:���%,���a 6���ly_X1�1� �Vs���&���[��?ѭH�:�:h'�&�'yQ�I�0����3.X?�����Ms�
����c�]��1�; �6�;��k����$���Y-ϵ�H˓�,/I?]���;O��͵��ˤtïV��K�6}�� g��Z����&NT[�$u6���t�b�̖��z=)x�g����E�R SS�����2�.���¨҇��5�I`�"���쓊�aK�:r���GԯT���$OSB�l�q{\�!���Ҝ�Z�<▭{K2¾36-e��t�Z?j�xJ�4ĸn�h��M�}�����dU���Y�Ij&�Ɗb�ܞT\(��pi��v�F˪���:O<�$��Y��e��)��{�S����'�`�׺!��&t�G�ҥ��������C  �C�~���͑�sB�p�Q��Iy�R"��:�]ۖ�ږng�~��a���|�_�s5��>B��+d��#��*X��Ⱥ���T�
y�s+HX�,�	rm0G��b��"���o)P��/�kߝ<dHl�'&��Ht{�� ��0B�[��(
��x� 7��$���ѹ/;�ʻS����׆���"^��D���Is	�x[.��l�7!��Q�7���l�_i��K��dQ���Gb�/6)�&�� %��"��O5&Q�n��������C=P]�/gy�O��oo�k��m8tss6�W�f�ӧZ5��x^�n���Q���OE��2�n�W��@�eA���,��o�U��yL��߰٢9�^I~�����Osl��)�d�
�P�;�{Ud\,��T.lg���-�3KJ��1�zUc��:�p��W�"7b�͝�抔hO�J��?��9`Y�����W�ˀ�>� �`��a�
���X��3^��Q�I�ء�0�["�m�
�[��Jf:���@4�|T�P+�z��[�a��5�Q��t�)���'�@��ݫy����6�^U� �����>I�1K�@�
�JR����a>�4u�J&�l�3��.���28R'�u�4�&�����p�����J��Q�N���#>�@��_4i.ȥ��L�R����`���ʈ�R��-����m[��}g�U/Ț��y[����=^�F�����G��eMp�*���iN���!�u'Q�Il�Z���mj��D�t���XJϔ_���"5�/�eH��T_셆y�ՠ��yM�
�iv�m�Ϛ���b1�X�I�"��ӇA1C����E�J�iV���G�٢��-��_+/fɞ�*1����۳��_�q
�t���ur��H�fy]ϰ������n,ё��ˊՀ�Z)7����dF����C��]Xn������Tw%���������͓ ����+M!��D�\.��Mf�?��F�����$ge?�,7B}8|���� �i��(J�=u���^�\�Ӥ������r�pA|t�*N��_}������^���$��Ê�����T���`Z�G�A���e@#�܁�H����EH��wo�xmP��9�%]��MŽVF�