LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE bchp_roots IS

type numarray IS ARRAY (0 TO 16383) OF integer;

constant negenum : numarray := (1,8737,13105,15289,16381,15839,15566,7783,11538,5769,10597,13971,14696,7348,3674,1837,
                   8631,13050,6525,11935,13678,6839,12154,6077,10751,14046,7023,12182,6091,10692,5346,
                   2673,10009,12717,15095,16218,8109,11767,13530,6765,12055,13738,6869,12107,13700,6850,
                   3425,9361,12393,14869,16171,15796,7898,3949,9623,12522,6261,11803,13612,6806,3403,
                   9348,4674,2337,9905,12665,15005,16239,15766,7883,11588,5794,2897,10121,12773,15059,
                   16200,8100,4050,2025,8661,13003,15172,7586,3793,9545,12421,14947,16144,8072,4036,
                   2018,1009,9177,13261,15303,16322,8161,11729,13513,14405,15875,15648,7824,3912,1956,
                   978,489,8917,13131,15236,7618,3809,9553,12425,14949,16147,15784,7892,3946,1973,
                   8699,13020,6510,3255,9338,4669,11071,14270,7135,12238,6119,10706,5353,10325,13835,
                   14628,7314,3657,9477,12451,14960,7480,3740,1870,935,9202,4601,10973,14159,14726,
                   7363,11328,5664,2832,1416,708,354,177,8825,13085,15279,16374,8187,11740,5870,
                   2935,10138,5069,11207,14274,7137,12241,13769,14533,15939,15616,7808,3904,1952,976,
                   488,244,122,61,8767,13118,6559,12014,6007,10650,5325,10311,13826,6913,12193,
                   13809,14553,15949,15623,15522,7761,11529,13477,14451,15896,7948,3974,1987,8640,4320,
                   2160,1080,540,270,135,8802,4401,10937,14205,14751,16110,8055,11674,5837,10567,
                   13954,6977,12161,13793,14545,15945,15621,15523,15472,7736,3868,1934,967,9154,4577,
                   10961,14153,14725,16099,15696,7848,3924,1962,981,9163,13252,6626,3313,9305,12301,
                   14887,16178,8089,11757,13527,14410,7205,11315,13368,6684,3342,1671,8546,4273,10873,
                   14109,14767,16118,8059,11676,5838,2919,10130,5065,11205,14275,14784,7392,3696,1848,
                   924,462,231,8786,4393,10933,14203,14748,7374,3687,9490,4745,11109,14227,14824,
                   7412,3706,1853,8639,13054,6527,11934,5967,10630,5315,10304,5152,2576,1288,644,
                   322,161,8817,13081,15277,16375,15834,7917,11607,13450,6725,12035,13728,6864,3432,
                   1716,858,429,8951,13146,6573,12023,13658,6829,12151,13722,6861,12103,13698,6849,
                   12097,13697,14561,15953,15625,15525,15475,15384,7692,3846,1923,8672,4336,2168,1084,
                   542,271,8870,4435,10888,5444,2722,1361,8329,12901,15123,16296,8148,4074,2037,
                   8667,13004,6502,3251,9336,4668,2334,1167,8294,4147,10808,5404,2702,1351,8322,
                   4161,10753,14113,14769,16121,15709,15503,15462,7731,11576,5788,2894,1447,8434,4217,
                   10781,14127,14774,7387,11340,5670,2835,10152,5076,2538,1269,8283,12812,6406,3203,
                   9312,4656,2328,1164,582,291,8880,4440,2220,1110,555,9012,4506,2253,9799,
                   12546,6273,11873,13585,14505,15989,15643,15532,7766,3883,9652,4826,2413,9879,12650,
                   6325,11899,13596,6798,3399,9346,4673,11009,14241,14833,16089,15693,15495,15458,7729,
                   11577,13501,14463,15902,7951,11686,5843,10568,5284,2642,1321,8373,12923,15132,7566,
                   3783,9538,4769,11121,14233,14829,16087,15690,7845,11635,13464,6732,3366,1683,8552,
                   4276,2138,1069,8247,12858,6429,11951,13686,6843,12156,6078,3039,10190,5095,11218,
                   5609,10453,13899,14596,7298,3649,9473,12449,14961,16153,15789,15607,15450,7725,11575,
                   13498,6749,12047,13734,6867,12104,6052,3026,1513,8405,12875,15108,7554,3777,9537,
                   12417,14945,16145,15785,15605,15451,15372,7686,3843,9632,4816,2408,1204,602,301,
                   8887,13178,6589,12031,13662,6831,12150,6075,10748,5374,2687,10014,5007,11238,5619,
                   10456,5228,2614,1307,8364,4182,2091,9780,4890,2445,9959,12626,6313,11893,13595,
                   14508,7254,3627,9524,4762,2381,9863,12642,6321,11897,13597,14511,15990,7995,11708,
                   5854,2927,10134,5067,11204,5602,2801,10073,12685,15079,16210,8105,11765,13531,14412,
                   7206,3603,9512,4756,2378,1189,8307,12824,6412,3206,1603,8448,4224,2112,1056,
                   528,264,132,66,33,8753,13113,15293,16383,15838,7919,11606,5803,10612,5306,
                   2653,9999,12710,6355,11848,5924,2962,1481,8389,12867,15104,7552,3776,1888,944,
                   472,236,118,59,8764,4382,2191,9830,4915,11192,5596,2798,1399,8346,4173,
                   10759,14114,7057,12265,13781,14539,15940,7970,3985,9705,12501,14923,16132,8066,4033,
                   9665,12481,14913,16129,15777,15601,15449,15373,15399,15410,7705,11565,13495,14458,7229,
                   11327,13374,6687,12078,6039,10730,5365,10331,13836,6918,3459,9440,4720,2360,1180,
                   590,295,8882,4441,10893,14183,14738,7369,11333,13315,14368,7184,3592,1796,898,
                   449,8897,13121,15233,16353,15825,15561,15429,15363,15392,7696,3848,1924,962,481,
                   8913,13129,15237,16355,15824,7912,3956,1978,989,9167,13254,6627,11984,5992,2996,
                   1498,749,9047,13194,6597,11971,13632,6816,3408,1704,852,426,213,8779,13060,
                   6530,3265,9281,12289,14881,16177,15801,15613,15455,15374,7687,11554,5777,10601,13973,
                   14699,16020,8010,4005,9715,12504,6252,3126,1563,8492,4246,2123,9732,4866,2433,
                   9953,12625,14985,16229,15763,15592,7796,3898,1949,8687,13014,6507,11924,5962,2981,
                   10227,12760,6380,3190,1595,8508,4254,2127,9734,4867,11168,5584,2792,1396,698,
                   349,8847,13158,6579,12024,6012,3006,1503,8398,4199,10770,5385,10405,13939,14616,
                   7308,3654,1827,8624,4312,2156,1078,539,9004,4502,2251,9796,4898,2449,9961,
                   12629,14987,16228,8114,4057,9677,12487,14914,7457,11441,13433,14365,15919,15670,7835,
                   11628,5814,2907,10124,5062,2531,9936,4968,2484,1242,621,8983,13226,6613,11979,
                   13636,6818,3409,9353,12389,14867,16168,8084,4042,2021,8659,13000,6500,3250,1625,
                   8461,12967,15218,7609,11517,13407,14350,7175,11298,5649,10537,14005,14715,16028,8014,
                   4007,9714,4857,11101,14223,14822,7411,11352,5676,2838,1419,8420,4210,2105,9789,
                   12607,15038,7519,11406,5703,10498,5249,10337,13841,14633,16053,15739,15516,7758,3879,
                   9650,4825,11085,14215,14818,7409,11353,13325,14375,15922,7961,11693,13559,14426,7213,
                   11319,13370,6685,12079,13750,6875,12108,6054,3027,10184,5092,2546,1273,8285,12815,
                   15142,7571,11496,5748,2874,1437,8431,12886,6443,11956,5978,2989,10231,12762,6381,
                   11863,13578,6789,12131,13712,6856,3428,1714,857,9101,13287,15314,7657,11477,13387,
                   14340,7170,3585,9505,12465,14969,16157,15791,15606,7803,11548,5774,2887,10114,5057,
                   11201,14273,14785,16065,15681,15489,15457,15377,15401,15413,15419,15420,7710,3855,9638,
                   4819,11080,5540,2770,1385,8341,12907,15124,7562,3781,9539,12416,6208,3104,1552,
                   776,388,194,97,8721,13097,15285,16379,15836,7918,3959,9626,4813,11079,14210,
                   7105,12225,13761,14529,15937,15617,15521,15473,15385,15405,15415,15418,7709,11567,13494,
                   6747,12044,6022,3011,10176,5088,2544,1272,636,318,159,8814,4407,10938,5469,
                   10383,13926,6963,12216,6108,3054,1527,8410,4205,10775,14122,7061,12267,13780,6890,
                   3445,9371,12396,6198,3099,9260,4630,2315,9892,4946,2473,9973,12635,14988,7494,
                   3747,9584,4792,2396,1198,599,8970,4485,10979,14160,7080,3540,1770,885,9115,
                   13292,6646,3323,9308,4654,2327,9898,4949,11147,14308,7154,3577,9437,12367,14854,
                   7427,11424,5712,2856,1428,714,357,8851,13160,6580,3290,1645,8471,12970,6485,
                   11915,13668,6834,3417,9357,12391,14866,7433,11429,13427,14360,7180,3590,1795,8608,
                   4304,2152,1076,538,269,8871,13170,6585,12029,13663,14478,7239,11266,5633,10529,
                   14001,14713,16029,15727,15510,7755,11524,5762,2881,10113,12769,15057,16201,15749,15587,
                   15440,7720,3860,1930,965,9155,13248,6624,3312,1656,828,414,207,8774,4387,
                   10928,5464,2732,1366,683,9076,4538,2269,9807,12550,6275,11872,5936,2968,1484,
                   742,371,8856,4428,2214,1107,8200,4100,2050,1025,8225,12849,15161,16317,15871,
                   15582,7791,11542,5771,10596,5298,2649,9997,12711,15090,7545,11421,13423,14358,7179,
                   11300,5650,2825,10149,12787,15064,7532,3766,1883,8588,4294,2147,9744,4872,2436,
                   1218,609,8977,13225,15349,16347,15820,7910,3955,9624,4812,2406,1203,8312,4156,
                   2078,1039,8230,4115,10792,5396,2698,1349,8323,12896,6448,3224,1612,806,403,
                   8936,4468,2234,1117,8207,12838,6419,11944,5972,2986,1493,8395,12868,6434,3217,
                   9321,12309,14891,16180,8090,4045,9671,12482,6241,11793,13609,14517,15995,15644,7822,
                   3911,9602,4801,11073,14209,14817,16081,15689,15493,15459,15376,7688,3844,1922,961,
                   9153,13249,15297,16321,15809,15553,15425,15361,15393,15409,15417,15421,15423,15422,7711,
                   11566,5783,10602,5301,10363,13852,6926,3463,9442,4721,11033,14253,14839,16090,8045,
                   11671,13546,6773,12059,13740,6870,3435,9364,4682,2341,9907,12664,6332,3166,1583,
                   8502,4251,10860,5430,2715,10092,5046,2523,9932,4966,2483,9976,4988,2494,1247,
                   8270,4135,10802,5401,10413,13943,14618,7309,11367,13330,6665,12069,13747,14584,7292,
                   3646,1823,8622,4311,10826,5413,10419,13944,6972,3486,1743,8518,4259,10864,5432,
                   2716,1358,679,9074,4537,11005,14175,14734,7367,11330,5665,10545,14009,14717,16031,
                   15726,7863,11642,5821,10623,13982,6991,12166,6083,10688,5344,2672,1336,668,334,
                   167,8818,4409,10941,14207,14750,7375,11334,5667,10544,5272,2636,1318,659,9064,
                   4532,2266,1133,8215,12842,6421,11947,13684,6842,3421,9359,12390,6195,11832,5916,
                   2958,1479,8386,4193,10769,14121,14773,16123,15708,7854,3927,9610,4805,11075,14208,
                   7104,3552,1776,888,444,222,111,8726,4363,10916,5458,2729,10101,12699,15084,
                   7542,3771,9596,4798,2399,9870,4935,11138,5569,10433,13889,14593,16033,15729,15513,
                   15469,15383,15402,7701,11563,13492,6746,3373,9399,12410,6205,11839,13630,6815,12142,
                   6071,10746,5373,10335,13838,6919,12194,6097,10697,14021,14659,16000,8000,4000,2000,
                   1000,500,250,125,8735,13102,6551,12010,6005,10651,14060,7030,3515,9468,4734,
                   2367,9918,4959,11150,5575,10434,5217,10257,13865,14645,16059,15740,7870,3935,9614,
                   4807,11074,5537,10481,13913,14605,16039,15730,7865,11645,13471,14446,7223,11322,5661,
                   10543,14006,7003,12172,6086,3043,10192,5096,2548,1274,637,8991,13230,6615,11978,
                   5989,10643,14056,7028,3514,1757,8527,12934,6467,11904,5952,2976,1488,744,372,
                   186,93,8719,13094,6547,12008,6004,3002,1501,8399,12870,6435,11952,5976,2988,
                   1494,747,9044,4522,2261,9803,12548,6274,3137,9217,12321,14897,16185,15805,15615,
                   15454,7727,11574,5787,10604,5302,2651,9996,4998,2499,9920,4960,2480,1240,620,
                   310,155,8812,4406,2203,9836,4918,2459,9964,4982,2491,9980,4990,2495,9982,
                   4991,11166,5583,10438,5219,10256,5128,2564,1282,641,9057,13201,15337,16341,15819,
                   15556,7778,3889,9657,12541,14943,16142,8071,11746,5873,10585,13965,14695,16018,8009,
                   11653,13539,14416,7208,3604,1802,901,9187,13264,6632,3316,1658,829,9151,13310,
                   6655,11998,5999,10646,5323,10308,5154,2577,10025,12725,15099,16220,8110,4055,9674,
                   4837,11091,14216,7108,3554,1777,8537,12941,15207,16274,8137,11717,13507,14400,7200,
                   3600,1800,900,450,225,8785,13065,15269,16371,15832,7916,3958,1979,8700,4350,
                   2175,9758,4879,11174,5587,10440,5220,2610,1305,8365,12919,15130,7565,11495,13394,
                   6697,12085,13755,14588,7294,3647,9534,4767,11118,5559,10490,5245,10271,13870,6935,
                   12202,6101,10699,14020,7010,3505,9465,12381,14863,16166,8083,11752,5876,2938,1469,
                   8447,12894,6447,11958,5979,10636,5318,2659,10000,5000,2500,1250,625,8985,13229,
                   15351,16346,8173,11735,13514,6757,12051,13736,6868,3434,1717,8571,12956,6478,3239,
                   9330,4665,11069,14271,14846,7423,11358,5679,10550,5275,10348,5174,2587,10028,5014,
                   2507,9924,4962,2481,9977,12637,14991,16230,8115,11768,5884,2942,1471,8446,4223,
                   10782,5391,10406,5203,10248,5124,2562,1281,8353,12913,15129,16301,15863,15578,7789,
                   11543,13482,6741,12043,13732,6866,3433,9365,12395,14868,7434,3717,9571,12432,6216,
                   3108,1554,777,9125,13299,15320,7660,3830,1915,8604,4302,2151,9746,4873,11173,
                   14323,14808,7404,3702,1851,8636,4318,2159,9750,4875,11172,5586,2793,10069,12683,
                   15076,7538,3769,9597,12447,14958,7479,11450,5725,10511,13990,6995,12168,6084,3042,
                   1521,8409,12877,15111,16290,8145,11721,13509,14403,15872,7936,3968,1984,992,496,
                   248,124,62,31,8750,4375,10922,5461,10379,13924,6962,3481,9453,12375,14858,
                   7429,11427,13424,6712,3356,1678,839,9090,4545,10945,14145,14721,16097,15697,15497,
                   15461,15379,15400,7700,3850,1925,8675,13008,6504,3252,1626,813,9143,13306,6653,
                   11999,13646,6823,12146,6073,10749,14047,14670,7335,11378,5689,10557,14015,14718,7359,
                   11390,5695,10558,5279,10350,5175,10298,5149,10287,13878,6939,12204,6102,3051,10196,
                   5098,2549,9947,12620,6310,3155,9224,4612,2306,1153,8289,12817,15145,16309,15867,
                   15580,7790,3895,9658,4829,11087,14214,7107,12224,6112,3056,1528,764,382,191,
                   8830,4415,10942,5471,10382,5191,10242,5121,10273,13873,14649,16061,15743,15518,7759,
                   11526,5763,10592,5296,2648,1324,662,331,8836,4418,2209,9841,12569,15021,16247,
                   15770,7885,11591,13442,6721,12033,13729,14577,15961,15629,15527,15474,7737,11581,13503,
                   14462,7231,11326,5663,10542,5271,10346,5173,10299,13884,6942,3471,9446,4723,11032,
                   5516,2758,1379,8336,4168,2084,1042,521,8997,13235,15352,7676,3838,1919,8606,
                   4303,10822,5411,10416,5208,2604,1302,651,9060,4530,2265,9805,12551,15010,7505,
                   11401,13413,14355,15912,7956,3978,1989,8643,12992,6496,3248,1624,812,406,203,
                   8772,4386,2193,9833,12565,15019,16244,8122,4061,9679,12486,6243,11792,5896,2948,
                   1474,737,9041,13193,15333,16339,15816,7908,3954,1977,8701,13023,15182,7591,11506,
                   5753,10525,13999,14710,7355,11388,5694,2847,10158,5079,11210,5605,10451,13896,6948,
                   3474,1737,8517,12931,15200,7600,3800,1900,950,475,8908,4454,2227,9848,4924,
                   2462,1231,8262,4131,10800,5400,2700,1350,675,9072,4536,2268,1134,567,9018,
                   4509,10991,14166,7083,12276,6138,3069,10207,12750,6375,11858,5929,10677,14075,14684,
                   7342,3671,9482,4741,11107,14224,7112,3556,1778,889,9117,13295,15318,7659,11476,
                   5738,2869,10171,12796,6398,3199,9246,4623,11046,5523,10472,5236,2618,1309,8367,
                   12918,6459,11964,5982,2991,10230,5115,11228,5614,2807,10074,5037,11255,14298,7149,
                   12247,13770,6885,12115,13704,6852,3426,1713,8569,12957,15215,16278,8139,11716,5858,
                   2929,10137,12781,15063,16202,8101,11763,13528,6764,3382,1691,8556,4278,2139,9740,
                   4870,2435,9952,4976,2488,1244,622,311,8890,4445,10895,14182,7091,12280,6140,
                   3070,1535,8414,4207,10774,5387,10404,5202,2601,10037,12731,15100,7550,3775,9598,
                   4799,11134,5567,10494,5247,10270,5135,10278,5139,10280,5140,2570,1285,8355,12912,
                   6456,3228,1614,807,9138,4569,10957,14151,14722,7361,11329,13313,14369,15921,15673,
                   15549,15487,15390,7695,11558,5779,10600,5300,2650,1325,8375,12922,6461,11967,13694,
                   6847,12158,6079,10750,5375,10334,5167,10294,5147,10284,5142,2571,10020,5010,2505,
                   9925,12611,14976,7488,3744,1872,936,468,234,117,8731,13100,6550,3275,9284,
                   4642,2321,9897,12661,15003,16236,8118,4059,9676,4838,2419,9880,4940,2470,1235,
                   8264,4132,2066,1033,8229,12851,15160,7580,3790,1895,8594,4297,10821,14083,14752,
                   7376,3688,1844,922,461,8903,13122,6561,12017,13657,14477,15975,15634,7817,11621,
                   13459,14440,7220,3610,1805,8615,13042,6521,11933,13679,14486,7243,11268,5634,2817,
                   10145,12785,15065,16205,15751,15586,7793,11545,13485,14455,15898,7949,11687,13554,6777,
                   12061,13743,14582,7291,11292,5646,2823,10146,5073,11209,14277,14787,16064,8032,4016,
                   2008,1004,502,251,8796,4398,2199,9834,4917,11195,14332,7166,3583,9438,4719,
                   11030,5515,10468,5234,2617,10045,12735,15102,7551,11422,5711,10502,5251,10336,5168,
                   2584,1292,646,323,8832,4416,2208,1104,552,276,138,69,8707,13088,6544,
                   3272,1636,818,409,8941,13143,15242,7621,11459,13376,6688,3344,1672,836,418,
                   209,8777,13061,15267,16368,8184,4092,2046,1023,9182,4591,10966,5483,10388,5194,
                   2597,10035,12728,6364,3182,1591,8506,4253,10863,14102,7051,12260,6130,3065,10205,
                   12751,15046,7523,11408,5704,2852,1426,713,9029,13187,15328,7664,3832,1916,958,
                   479,8910,4455,10898,5449,10373,13923,14608,7304,3652,1826,913,9193,13269,15307,
                   16324,8162,4081,9689,12493,14919,16130,8065,11745,13521,14409,15877,15651,15536,7768,
                   3884,1942,971,9156,4578,2289,9817,12557,15015,16242,8121,11773,13535,14414,7207,
                   11314,5657,10541,14007,14714,7357,11391,13342,6671,12070,6035,10728,5364,2682,1341,
                   8383,12926,6463,11966,5983,10638,5319,10306,5153,10289,13881,14653,16063,15742,7871,
                   11646,5823,10622,5311,10366,5183,10302,5151,10286,5143,10282,5141,10283,13876,6938,
                   3469,9447,12370,6185,11829,13627,14524,7262,3631,9526,4763,11116,5558,2779,10060,
                   5030,2515,9928,4964,2482,1241,8269,12807,15138,7569,11497,13397,14347,15908,7954,
                   3977,9701,12499,14920,7460,3730,1865,8581,13027,15184,7592,3796,1898,949,9211,
                   13276,6638,3319,9306,4653,11063,14266,7133,12239,13766,6883,12112,6056,3028,1514,
                   757,9051,13196,6598,3299,9296,4648,2324,1162,581,8963,13216,6608,3304,1652,
                   826,413,8943,13142,6571,12020,6010,3005,10239,12766,6383,11862,5931,10676,5338,
                   2669,10007,12714,6357,11851,13572,6786,3393,9345,12385,14865,16169,15797,15611,15452,
                   7726,3863,9642,4821,11083,14212,7106,3553,9425,12361,14853,16163,15792,7896,3948,
                   1974,987,9164,4582,2291,9816,4908,2454,1227,8260,4130,2065,9769,12597,15035,
                   16252,8126,4063,9678,4839,11090,5545,10485,13915,14604,7302,3651,9472,4736,2368,
                   1184,592,296,148,74,37,8755,13112,6556,3278,1639,8466,4233,10853,14099,
                   14760,7380,3690,1845,8635,13052,6526,3263,9342,4671,11070,5535,10478,5239,10266,
                   5133,10279,13874,6937,12205,13815,14554,7277,11287,13354,6677,12075,13748,6874,3437,
                   9367,12394,6197,11835,13628,6814,3407,9350,4675,11008,5504,2752,1376,688,344,
                   172,86,43,8756,4378,2189,9831,12562,6281,11877,13587,14504,7252,3626,1813,
                   8619,13044,6522,3261,9343,12318,6159,11814,5907,10664,5332,2666,1333,8379,12924,
                   6462,3231,9326,4663,11066,5533,10479,13910,6955,12212,6106,3053,10199,12746,6373,
                   11859,13576,6788,3394,1697,8561,12953,15213,16279,15850,7925,11611,13452,6726,3363,
                   9392,4696,2348,1174,587,8964,4482,2241,9793,12545,15009,16241,15769,15597,15447,
                   15370,7685,11555,13488,6744,3372,1686,843,9092,4546,2273,9809,12553,15013,16243,
                   15768,7884,3942,1971,8696,4348,2174,1087,8254,4127,10798,5399,10410,5205,10251,
                   13860,6930,3465,9445,12371,14856,7428,3714,1857,8577,13025,15185,16265,15845,15571,
                   15432,7716,3858,1929,8677,13011,15176,7588,3794,1897,8597,13035,15188,7594,3797,
                   9547,12420,6210,3105,9265,12345,14909,16191,15806,7903,11598,5799,10610,5305,10365,
                   13855,14638,7319,11370,5685,10555,14012,7006,3503,9462,4731,11036,5518,2759,10050,
                   5025,11249,14297,14797,16071,15682,7841,11633,13465,14445,15895,15658,7829,11627,13460,
                   6730,3365,9395,12408,6204,3102,1551,8486,4243,10856,5428,2714,1357,8327,12898,
                   6449,11961,13693,14495,15982,7991,11706,5853,10575,13958,6979,12160,6080,3040,1520,
                   760,380,190,95,8718,4359,10914,5457,10377,13925,14611,16040,8020,4010,2005,
                   8651,12996,6498,3249,9337,12317,14895,16182,8091,11756,5878,2939,10140,5070,2535,
                   9938,4969,11157,14315,14804,7402,3701,9499,12460,6230,3115,9268,4634,2317,9895,
                   12658,6329,11901,13599,14510,7255,11274,5637,10531,14000,7000,3500,1750,875,9108,
                   4554,2277,9811,12552,6276,3138,1569,8497,12985,15229,16287,15854,7927,11610,5805,
                   10615,13978,6989,12167,13794,6897,12121,13709,14567,15954,7977,11701,13563,14428,7214,
                   3607,9514,4757,11115,14228,7114,3557,9427,12360,6180,3090,1545,8485,12979,15224,
                   7612,3806,1903,8598,4299,10820,5410,2705,10089,12693,15083,16212,8106,4053,9675,
                   12484,6242,3121,9273,12349,14911,16190,8095,11758,5879,10586,5293,10359,13850,6925,
                   12199,13810,6905,12125,13711,14566,7283,11288,5644,2822,1411,8416,4208,2104,1052,
                   526,263,8866,4433,10889,14181,14739,16104,8052,4026,2013,8655,12998,6499,11920,
                   5960,2980,1490,745,9045,13195,15332,7666,3833,9565,12431,14950,7475,11448,5724,
                   2862,1431,8426,4213,10779,14124,7062,3531,9412,4706,2353,9913,12669,15007,16238,
                   8119,11770,5885,10591,13966,6983,12162,6081,10689,14017,14657,16001,15713,15505,15465,
                   15381,15403,15412,7706,3853,9639,12530,6265,11805,13615,14518,7259,11276,5638,2819,
                   10144,5072,2536,1268,634,317,8895,13182,6591,12030,6015,10654,5327,10310,5155,
                   10288,5144,2572,1286,643,9056,4528,2264,1132,566,283,8876,4438,2219,9844,
                   4922,2461,9967,12630,6315,11892,5946,2973,10223,12758,6379,11860,5930,2965,10219,
                   12756,6378,3189,9243,12332,6166,3083,9252,4626,2313,9893,12659,15000,7500,3750,
                   1875,8584,4292,2146,1073,8249,12861,15167,16318,8159,11726,5863,10578,5289,10357,
                   13851,14636,7318,3659,9476,4738,2369,9857,12641,14993,16233,15765,15595,15444,7722,
                   3861,9643,12532,6266,3133,9279,12350,6175,11822,5911,10666,5333,10315,13828,6914,
                   3457,9441,12369,14857,16165,15795,15608,7804,3902,1951,8686,4343,10842,5421,10423,
                   13946,6973,12223,13822,6911,12126,6063,10742,5371,10332,5166,2583,10026,5013,11243,
                   14292,7146,3573,9435,12364,6182,3091,9256,4628,2314,1157,8291,12816,6408,3204,
                   1602,801,9137,13305,15325,16335,15814,7907,11600,5800,2900,1450,725,9035,13188,
                   6594,3297,9297,12297,14885,16179,15800,7900,3950,1975,8698,4349,10847,14094,7047,
                   12258,6129,10713,14029,14663,16002,8001,11649,13537,14417,15881,15653,15539,15480,7740,
                   3870,1935,8678,4339,10840,5420,2710,1355,8324,4162,2081,9777,12601,15037,16255,
                   15774,7887,11590,5795,10608,5304,2652,1326,663,9066,4533,11003,14172,7086,3543,
                   9418,4709,11027,14248,7124,3562,1781,8539,12940,6470,3235,9328,4664,2332,1166,
                   583,8962,4481,10977,14161,14729,16101,15699,15496,7748,3874,1937,8681,13013,15179,
                   16260,8130,4065,9681,12489,14917,16131,15776,7888,3944,1972,986,493,8919,13130,
                   6565,12019,13656,6828,3414,1707,8564,4282,2141,9743,12582,6291,11880,5940,2970,
                   1485,8391,12866,6433,11953,13689,14493,15983,15638,7819,11620,5810,2905,10125,12775,
                   15058,7529,11413,13419,14356,7178,3589,9507,12464,6232,3116,1558,779,9124,4562,
                   2281,9813,12555,15012,7506,3753,9589,12443,14956,7478,3739,9580,4790,2395,9868,
                   4934,2467,9968,4984,2492,1246,623,8982,4491,10980,5490,2745,10109,12703,15086,
                   7543,11418,5709,10503,13986,6993,12169,13797,14547,15944,7972,3986,1993,8645,12995,
                   15168,7584,3792,1896,948,474,237,8791,13066,6533,12003,13648,6824,3412,1706,
                   853,9099,13284,6642,3321,9309,12303,14886,7443,11432,5716,2858,1429,8427,12884,
                   6442,3221,9323,12308,6154,3077,9251,12336,6168,3084,1542,771,9120,4560,2280,
                   1140,570,285,8879,13174,6587,12028,6014,3007,10238,5119,11230,5615,10454,5227,
                   10260,5130,2565,10019,12720,6360,3180,1590,795,9132,4566,2283,9812,4906,2453,
                   9963,12628,6314,3157,9227,12324,6162,3081,9253,12339,14904,7452,3726,1863,8578,
                   4289,10817,14081,14753,16113,15705,15501,15463,15378,7689,11557,13491,14456,7228,3614,
                   1807,8614,4307,10824,5412,2706,1353,8325,12899,15120,7560,3780,1890,945,9209,
                   13277,15311,16326,8163,11728,5864,2932,1466,733,9039,13190,6595,11968,5984,2992,
                   1496,748,374,187,8828,4414,2207,9838,4919,11194,5597,10447,13894,6947,12208,
                   6104,3052,1526,763,9052,4526,2263,9802,4901,11187,14328,7164,3582,1791,8542,
                   4271,10870,5435,10428,5214,2607,10038,5019,11244,5622,2811,10076,5038,2519,9930,
                   4965,11155,14312,7156,3578,1789,8543,12942,6471,11906,5953,10625,14049,14673,16009,
                   15717,15507,15464,7732,3866,1933,8679,13010,6505,11925,13675,14484,7242,3621,9523,
                   12472,6236,3118,1559,8490,4245,10859,14100,7050,3525,9411,12352,6176,3088,1544,
                   772,386,193,8769,13057,15265,16369,15833,15565,15431,15362,7681,11553,13489,14457,
                   15901,15663,15542,7771,11532,5766,2883,10112,5056,2528,1264,632,316,158,79,
                   8710,4355,10912,5456,2728,1364,682,341,8843,13156,6578,3289,9293,12295,14882,
                   7441,11433,13429,14363,15916,7958,3979,9700,4850,2425,9885,12655,14998,7499,11396,
                   5698,2849,10161,12793,15069,16207,15750,7875,11584,5792,2896,1448,724,362,181,
                   8827,13084,6542,3271,9282,4641,11057,14265,14845,16095,15694,7847,11634,5817,10621,
                   13983,14702,7351,11386,5693,10559,14014,7007,12174,6087,10690,5345,10321,13833,14629,
                   16051,15736,7868,3934,1967,8694,4347,10844,5422,2711,10090,5045,11259,14300,7150,
                   3575,9434,4717,11031,14250,7125,12235,13764,6882,3441,9369,12397,14871,16170,8085,
                   11755,13524,6762,3381,9403,12412,6206,3103,9262,4631,11050,5525,10475,13908,6954,
                   3477,9451,12372,6186,3093,9259,12340,6170,3085,9255,12338,6169,11821,13623,14522,
                   7261,11279,13350,6675,12072,6036,3018,1509,8403,12872,6436,3218,1609,8453,12963,
                   15216,7608,3804,1902,951,9210,4605,10975,14158,7079,12274,6137,10717,14031,14662,
                   7331,11376,5688,2844,1422,711,9026,4513,10993,14169,14733,16103,15698,7849,11637,
                   13467,14444,7222,3611,9516,4758,2379,9860,4930,2465,9969,12633,14989,16231,15762,
                   7881,11589,13443,14432,7216,3608,1804,902,451,8896,4448,2224,1112,556,278,
                   139,8804,4402,2201,9837,12567,15018,7509,11403,13412,6706,3353,9389,12407,14874,
                   7437,11431,13426,6713,12093,13759,14590,7295,11294,5647,10534,5267,10344,5172,2586,
                   1293,8359,12914,6457,11965,13695,14494,7247,11270,5635,10528,5264,2632,1316,658,
                   329,8837,13155,15248,7624,3812,1906,953,9213,13279,15310,7655,11474,5737,10517,
                   13995,14708,7354,3677,9487,12454,6227,11784,5892,2946,1473,8385,12865,15105,16289,
                   15857,15577,15437,15367,15394,7697,11561,13493,14459,15900,7950,3975,9698,4849,11097,
                   14221,14823,16082,8041,11669,13547,14420,7210,3605,9515,12468,6234,3117,9271,12346,
                   6173,11823,13622,6811,12140,6070,3035,10188,5094,2547,9944,4972,2486,1243,8268,
                   4134,2067,9768,4884,2442,1221,8259,12800,6400,3200,1600,800,400,200,100,
                   50,25,8749,13111,15290,7645,11471,13382,6691,12080,6040,3020,1510,755,9048,
                   4524,2262,1131,8212,4106,2053,9763,12592,6296,3148,1574,787,9128,4564,2282,
                   1141,8219,12844,6422,3211,9316,4658,2329,9901,12663,15002,7501,11399,13410,6705,
                   12089,13757,14591,15966,7983,11702,5851,10572,5286,2643,9992,4996,2498,1249,8273,
                   12809,15141,16307,15864,7932,3966,1983,8702,4351,10846,5423,10422,5211,10252,5126,
                   2563,10016,5008,2504,1252,626,313,8893,13183,15262,7631,11462,5731,10512,5256,
                   2628,1314,657,9065,13205,15339,16340,8170,4085,9691,12492,6246,3123,9272,4636,
                   2318,1159,8290,4145,10809,14141,14783,16126,8063,11678,5839,10566,5283,10352,5176,
                   2588,1294,647,9058,4529,11001,14173,14735,16102,8051,11672,5836,2918,1459,8440,
                   4220,2110,1055,8238,4119,10794,5397,10411,13940,6970,3485,9455,12374,6187,11828,
                   5914,2957,10215,12754,6377,11861,13579,14500,7250,3625,9525,12475,14972,7486,3743,
                   9582,4791,11130,5565,10495,13918,6959,12214,6107,10700,5350,2675,10008,5004,2502,
                   1251,8272,4136,2068,1034,517,8995,13232,6616,3308,1654,827,9148,4574,2287,
                   9814,4907,11188,5594,2797,10071,12682,6341,11843,13568,6784,3392,1696,848,424,
                   212,106,53,8763,13116,6558,3279,9286,4643,11056,5528,2764,1382,691,9080,
                   4540,2270,1135,8214,4107,10788,5394,2697,10085,12691,15080,7540,3770,1885,8591,
                   13030,6515,11928,5964,2982,1491,8392,4196,2098,1049,8237,12855,15162,7581,11503,
                   13398,6699,12084,6042,3021,10183,12738,6369,11857,13577,14501,15987,15640,7820,3910,
                   1955,8688,4344,2172,1086,543,9006,4503,10986,5493,10395,13932,6966,3483,9452,
                   4726,2363,9916,4958,2479,9974,4987,11164,5582,2791,10066,5033,11253,14299,14796,
                   7398,3699,9496,4748,2374,1187,8304,4152,2076,1038,519,8994,4497,10985,14165,
                   14731,16100,8050,4025,9725,12511,14926,7463,11442,5721,10509,13991,14706,7353,11389,
                   13343,14382,7191,11306,5653,10539,14004,7002,3501,9463,12378,6189,11831,13626,6813,
                   12143,13718,6859,12100,6050,3025,10185,12741,15043,16192,8096,4048,2024,1012,506,
                   253,8799,13070,6535,12002,6001,10649,14061,14679,16010,8005,11651,13536,6768,3384,
                   1692,846,423,8946,4473,10909,14191,14742,7371,11332,5666,2833,10153,12789,15067,
                   16204,8102,4051,9672,4836,2418,1209,8317,12831,15150,7575,11498,5749,10523,13996,
                   6998,3499,9460,4730,2365,9919,12670,6335,11902,5951,10686,5343,10318,5159,10290,
                   5145,10285,13879,14650,7325,11375,13334,6667,12068,6034,3017,10181,12739,15040,7520,
                   3760,1880,940,470,235,8788,4394,2197,9835,12564,6282,3141,9219,12320,6160,
                   3080,1540,770,385,8929,13137,15241,16357,15827,15560,7780,3890,1945,8685,13015,
                   15178,7589,11507,13400,6700,3350,1675,8548,4274,2137,9741,12583,15026,7513,11405,
                   13415,14354,7177,11301,13363,14392,7196,3598,1799,8610,4305,10825,14085,14755,16112,
                   8056,4028,2014,1007,9174,4587,10964,5482,2741,10107,12700,6350,3175,9234,4617,
                   11045,14259,14840,7420,3710,1855,8638,4319,10830,5415,10418,5209,10253,13863,14642,
                   7321,11373,13335,14378,7189,11307,13364,6682,3341,9383,12402,6201,11837,13631,14526,
                   7263,11278,5639,10530,5265,10345,13845,14635,16052,8026,4013,9719,12506,6253,11799,
                   13610,6805,12139,13716,6858,3429,9363,12392,6196,3098,1549,8487,12978,6489,11917,
                   13671,14482,7241,11269,13347,14384,7192,3596,1798,899,9184,4592,2296,1148,574,
                   287,8878,4439,10890,5445,10371,13920,6960,3480,1740,870,435,8952,4476,2238,
                   1119,8206,4103,10786,5393,10409,13941,14619,16044,8022,4011,9716,4858,2429,9887,
                   12654,6327,11898,5949,10687,14078,7039,12190,6095,10694,5347,10320,5160,2580,1290,
                   645,9059,13200,6600,3300,1650,825,9149,13311,15326,7663,11478,5739,10516,5258,
                   2629,9987,12704,6352,3176,1588,794,397,8935,13138,6569,12021,13659,14476,7238,
                   3619,9520,4760,2380,1190,595,8968,4484,2242,1121,8209,12841,15157,16315,15868,
                   7934,3967,9630,4815,11078,5539,10480,5240,2620,1310,655,9062,4531,11000,5500,
                   2750,1375,8334,4167,10754,5377,10401,13937,14617,16045,15735,15514,7757,11527,13474,
                   6737,12041,13733,14579,15960,7980,3990,1995,8644,4322,2161,9753,12589,15031,16250,
                   8125,11775,13534,6767,12054,6027,10724,5362,2681,10013,12719,15094,7547,11420,5710,
                   2855,10162,5081,11213,14279,14786,7393,11345,13321,14373,15923,15672,7836,3918,1959,
                   8690,4345,10845,14095,14758,7379,11336,5668,2834,1417,8421,12883,15112,7556,3778,
                   1889,8593,13033,15189,16267,15844,7922,3961,9629,12527,14934,7467,11444,5722,2861,
                   10167,12794,6397,11871,13582,6791,12130,6065,10745,14045,14671,16006,8003,11648,5824,
                   2912,1456,728,364,182,91,8716,4358,2179,9824,4912,2456,1228,614,307,
                   8888,4444,2222,1111,8202,4101,10787,14128,7064,3532,1766,883,9112,4556,2278,
                   1139,8216,4108,2054,1027,8224,4112,2056,1028,514,257,8865,13169,15257,16365,
                   15831,15562,7781,11539,13480,6740,3370,1685,8555,12948,6474,3237,9331,12312,6156,
                   3078,1539,8480,4240,2120,1060,530,265,8869,13171,15256,7628,3814,1907,8600,
                   4300,2150,1075,8248,4124,2062,1031,8226,4113,10793,14133,14779,16124,8062,4031,
                   9726,4863,11102,5551,10486,5243,10268,5134,2567,10018,5009,11241,14293,14795,16068,
                   8034,4017,9721,12509,14927,16134,8067,11744,5872,2936,1468,734,367,8854,4427,
                   10884,5442,2721,10097,12697,15085,16215,15754,7877,11587,13440,6720,3360,1680,840,
                   420,210,105,8725,13099,15284,7642,3821,9559,12426,6213,11779,13600,6800,3400,
                   1700,850,425,8949,13147,15244,7622,3811,9552,4776,2388,1194,597,8971,13220,
                   6610,3305,9301,12299,14884,7442,3721,9573,12435,14952,7476,3738,1869,8583,13026,
                   6513,11929,13677,14487,15978,7989,11707,13564,6782,3391,9406,4703,11022,5511,10466,
                   5233,10265,13869,14647,16058,8029,11663,13542,6771,12056,6028,3014,1507,8400,4200,
                   2100,1050,525,8999,13234,6617,11981,13639,14466,7233,11265,13345,14385,15929,15677,
                   15551,15486,7743,11582,5791,10606,5303,10362,5181,10303,13886,6943,12206,6103,10698,
                   5349,10323,13832,6916,3458,1729,8513,12929,15201,16273,15849,15573,15435,15364,7682,
                   3841,9633,12529,14937,16141,15783,15602,7801,11549,13487,14454,7227,11324,5662,2831,
                   10150,5075,11208,5604,2802,1401,8349,12911,15126,7563,11492,5746,2873,10173,12799,
                   15070,7535,11414,5707,10500,5250,2625,9985,12705,15089,16217,15757,15591,15442,7721,
                   11573,13499,14460,7230,3615,9518,4759,11114,5557,10491,13916,6958,3479,9450,4725,
                   11035,14252,7126,3563,9428,4714,2357,9915,12668,6334,3167,9230,4615,11042,5521,
                   10473,13909,14603,16036,8018,4009,9717,12507,14924,7462,3731,9576,4788,2394,1197,
                   8311,12826,6413,11943,13682,6841,12157,13727,14574,7287,11290,5645,10535,14002,7001,
                   12173,13799,14546,7273,11285,13355,14388,7194,3597,9511,12466,6233,11789,13607,14514,
                   7257,11277,13351,14386,7193,11309,13367,14394,7197,11311,13366,6683,12076,6038,3019,
                   10180,5090,2545,9945,12621,14983,16226,8113,11769,13533,14415,15878,7939,11680,5840,
                   2920,1460,730,365,8855,13162,6581,12027,13660,6830,3415,9354,4677,11011,14240,
                   7120,3560,1780,890,445,8959,13150,6575,12022,6011,10652,5326,2663,10002,5001,
                   11237,14291,14792,7396,3698,1849,8637,13055,15198,7599,11510,5755,10524,5262,2631,
                   9986,4993,11233,14289,14793,16069,15683,15488,7744,3872,1936,968,484,242,121,
                   8733,13103,15286,7643,11468,5734,2867,10168,5084,2542,1271,8282,4141,10807,14138,
                   7069,12271,13782,6891,12116,6058,3029,10187,12740,6370,3185,9241,12333,14903,16186,
                   8093,11759,13526,6763,12052,6026,3013,10179,12736,6368,3184,1592,796,398,199,
                   8770,4385,10929,14201,14749,16111,15702,7851,11636,5818,2909,10127,12774,6387,11864,
                   5932,2966,1483,8388,4194,2097,9785,12605,15039,16254,8127,11774,5887,10590,5295,
                   10358,5179,10300,5150,2575,10022,5011,11240,5620,2810,1405,8351,12910,6455,11962,
                   5981,10639,14054,7027,12184,6092,3046,1523,8408,4204,2102,1051,8236,4118,2059,
                   9764,4882,2441,9957,12627,14984,7492,3746,1873,8585,13029,15187,16264,8132,4066,
                   2033,8665,13005,15175,16258,8129,11713,13505,14401,15873,15649,15537,15481,15389,15407,
                   15414,7707,11564,5782,2891,10116,5058,2529,9937,12617,14981,16227,15760,7880,3940,
                   1970,985,9165,13255,15298,7649,11473,13385,14341,15907,15664,7832,3916,1958,979,
                   9160,4580,2290,1145,8221,12847,15158,7579,11500,5750,2875,10172,5086,2543,9942,
                   4971,11156,5578,2789,10067,12680,6340,3170,1585,8505,12989,15231,16286,8143,11718,
                   5859,10576,5288,2644,1322,661,9067,13204,6602,3301,9299,12296,6148,3074,1537,
                   8481,12977,15225,16285,15855,15574,7787,11540,5770,2885,10115,12768,6384,3192,1596,
                   798,399,8934,4467,10904,5452,2726,1363,8328,4164,2082,1041,8233,12853,15163,
                   16316,8158,4079,9686,4843,11092,5546,2773,10059,12676,6338,3169,9233,12329,14901,
                   16187,15804,7902,3951,9622,4811,11076,5538,2769,10057,12677,15075,16208,8104,4052,
                   2026,1013,9179,13260,6630,3315,9304,4652,2326,1163,8292,4146,2073,9773,12599,
                   15034,7517,11407,13414,6707,12088,6044,3022,1511,8402,4201,10773,14123,14772,7386,
                   3693,9495,12458,6229,11787,13604,6802,3401,9349,12387,14864,7432,3716,1858,929,
                   9201,13273,15309,16327,15810,7905,11601,13449,14437,15891,15656,7828,3914,1957,8691,
                   13016,6508,3254,1627,8460,4230,2115,9728,4864,2432,1216,608,304,152,76,
                   38,19,8744,4372,2186,1093,8195,12832,6416,3208,1604,802,401,8937,13141,
                   15243,16356,8178,4089,9693,12495,14918,7459,11440,5720,2860,1430,715,9028,4514,
                   2257,9801,12549,15011,16240,8120,4060,2030,1015,9178,4589,10967,14154,7077,12275,
                   13784,6892,3446,1723,8572,4286,2143,9742,4871,11170,5585,10441,13893,14595,16032,
                   8016,4008,2004,1002,501,8923,13132,6566,3283,9288,4644,2322,1161,8293,12819,
                   15144,7572,3786,1893,8595,13032,6516,3258,1629,8463,12966,6483,11912,5956,2978,
                   1489,8393,12869,15107,16288,8144,4072,2036,1018,509,8927,13134,6567,12018,6009,
                   10653,14063,14678,7339,11380,5690,2845,10159,12790,6395,11868,5934,2967,10218,5109,
                   11227,14284,7142,3571,9432,4716,2358,1179,8300,4150,2075,9772,4886,2443,9956,
                   4978,2489,9981,12639,14990,7495,11394,5697,10497,13985,14705,16025,15725,15511,15466,
                   7733,11579,13500,6750,3375,9398,4699,11020,5510,2755,10048,5024,2512,1256,628,
                   314,157,8815,13078,6539,12004,6002,3001,10237,12767,15054,7527,11410,5705,10501,
                   13987,14704,7352,3676,1838,919,9194,4597,10971,14156,7078,3539,9416,4708,2354,
                   1177,8301,12823,15146,7573,11499,13396,6698,3349,9387,12404,6202,3101,9263,12342,
                   6171,11820,5910,2955,10212,5106,2553,9949,12623,14982,7491,11392,5696,2848,1424,
                   712,356,178,89,8717,13095,15282,7641,11469,13383,14338,7169,11297,13361,14393,
                   15933,15679,15550,7775,11534,5767,10594,5297,10361,13853,14639,16054,8027,11660,5830,
                   2915,10128,5064,2532,1266,633,8989,13231,15350,7675,11484,5742,2871,10170,5085,
                   11215,14278,7139,12240,6120,3060,1530,765,9055,13198,6599,11970,5985,10641,14057,
                   14677,16011,15716,7858,3929,9613,12519,14930,7465,11445,13435,14364,7182,3591,9506,
                   4753,11113,14229,14827,16084,8042,4021,9723,12508,6254,3127,9274,4637,11055,14262,
                   7131,12236,6118,3059,10200,5100,2550,1275,8284,4142,2071,9770,4885,11179,14324,
                   7162,3581,9439,12366,6183,11826,5913,10669,14071,14682,7341,11383,13338,6669,12071,
                   13746,6873,12109,13703,14562,7281,11289,13357,14391,15930,7965,11695,13558,6779,12060,
                   6030,3015,10178,5089,11217,14281,14789,16067,15680,7840,3920,1960,980,490,245,
                   8795,13068,6534,3267,9280,4640,2320,1160,580,290,145,8809,13077,15275,16372,
                   8186,4093,9695,12494,6247,11794,5897,10661,14067,14680,7340,3670,1835,8628,4314,
                   2157,9751,12586,6293,11883,13588,6794,3397,9347,12384,6192,3096,1548,774,387,
                   8928,4464,2232,1116,558,279,8874,4437,10891,14180,7090,3545,9421,12359,14850,
                   7425,11425,13425,14361,15917,15671,15546,7773,11535,13478,6739,12040,6020,3010,1505,
                   8401,12873,15109,16291,15856,7928,3964,1982,991,9166,4583,10962,5481,10389,13931,
                   14612,7306,3653,9475,12448,6224,3112,1556,778,389,8931,13136,6568,3284,1642,
                   821,9147,13308,6654,3327,9310,4655,11062,5531,10476,5238,2619,10044,5022,2511,
                   9926,4963,11152,5576,2788,1394,697,9085,13215,15342,7671,11482,5741,10519,13994,
                   6997,12171,13796,6898,3449,9373,12399,14870,7435,11428,5714,2857,10165,12795,15068,
                   7534,3767,9594,4797,11135,14238,7119,12230,6115,10704,5352,2676,1338,669,9071,
                   13206,6603,11972,5986,2993,10233,12765,15055,16198,8099,11760,5880,2940,1470,735,
                   9038,4519,10994,5497,10397,13935,14614,7307,11364,5682,2841,10157,12791,15066,7533,
                   11415,13418,6709,12091,13756,6878,3439,9366,4683,11012,5506,2753,10049,12673,15073,
                   16209,15753,15589,15443,15368,7684,3842,1921,8673,13009,15177,16261,15843,15568,7784,
                   3892,1946,973,9159,13250,6625,11985,13641,14469,15971,15632,7816,3908,1954,977,
                   9161,13253,15299,16320,8160,4080,2040,1020,510,255,8798,4399,10934,5467,10380,
                   5190,2595,10032,5016,2508,1254,627,8984,4492,2246,1123,8208,4104,2052,1026,
                   513,8993,13233,15353,16349,15823,15558,7779,11536,5768,2884,1442,721,9033,13189,
                   15331,16336,8168,4084,2042,1021,9183,13262,6631,11986,5993,10645,14059,14676,7338,
                   3669,9483,12452,6226,3113,9269,12347,14908,7454,3727,9574,4787,11128,5564,2782,
                   1391,8342,4171,10756,5378,2689,10081,12689,15081,16213,15755,15588,7794,3897,9661,
                   12543,14942,7471,11446,5723,10508,5254,2627,9984,4992,2496,1248,624,312,156,
                   78,39,8754,4377,10925,14199,14746,7373,11335,13314,6657,12065,13745,14585,15965,
                   15631,15526,7763,11528,5764,2882,1441,8433,12889,15117,16295,15858,7929,11613,13455,
                   14438,7219,11320,5660,2830,1415,8418,4209,10777,14125,14775,16122,8061,11679,13550,
                   6775,12058,6029,10727,14034,7017,12181,13803,14548,7274,3637,9531,12476,6238,3119,
                   9270,4635,11052,5526,2763,10052,5026,2513,9929,12613,14979,16224,8112,4056,2028,
                   1014,507,8924,4462,2231,9850,4925,11199,14334,7167,12254,6127,10710,5355,10324,
                   5162,2581,10027,12724,6362,3181,9239,12330,6165,11819,13620,6810,3405,9351,12386,
                   6193,11833,13629,14527,15998,7999,11710,5855,10574,5287,10354,5177,10301,13887,14654,
                   7327,11374,5687,10554,5277,10351,13846,6923,12196,6098,3049,10197,12747,15044,7522,
                   3761,9593,12445,14959,16150,8075,11748,5874,2937,10141,12783,15062,7531,11412,5706,
                   2853,10163,12792,6396,3198,1599,8510,4255,10862,5431,10426,5213,10255,13862,6931,
                   12200,6100,3050,1525,8411,12876,6438,3219,9320,4660,2330,1165,8295,12818,6409,
                   11941,13683,14488,7244,3622,1811,8616,4308,2154,1077,8251,12860,6430,3215,9318,
                   4659,11064,5532,2766,1383,8338,4169,10757,14115,14768,7384,3692,1846,923,9196,
                   4598,2299,9820,4910,2455,9962,4981,11163,14316,7158,3579,9436,4718,2359,9914,
                   4957,11151,14310,7155,12248,6124,3062,1531,8412,4206,2103,9786,4893,11183,14326,
                   7163,12252,6126,3063,10202,5101,11223,14282,7141,12243,13768,6884,3442,1721,8573,
                   12959,15214,7607,11514,5757,10527,13998,6999,12170,6085,10691,14016,7008,3504,1752,
                   876,438,219,8780,4390,2195,9832,4916,2458,1229,8263,12802,6401,11937,13681,
                   14489,15981,15639,15530,7765,11531,13476,6738,3369,9397,12411,14876,7438,3719,9570,
                   4785,11129,14237,14831,16086,8043,11668,5834,2917,10131,12776,6388,3194,1597,8511,
                   12990,6495,11918,5959,10626,5313,10305,13825,14625,16049,15737,15517,15471,15382,7691,
                   11556,5778,2889,10117,12771,15056,7528,3764,1882,941,9207,13274,6637,11991,13642,
                   6821,12147,13720,6860,3430,1715,8568,4284,2142,1071,8246,4123,10796,5398,2699,
                   10084,5042,2521,9933,12615,14978,7489,11393,13409,14353,15913,15669,15547,15484,7742,
                   3871,9646,4823,11082,5541,10483,13912,6956,3478,1739,8516,4258,2129,9737,12581,
                   15027,16248,8124,4062,2031,8662,4331,10836,5418,2709,10091,12692,6346,3173,9235,
                   12328,6164,3082,1541,8483,12976,6488,3244,1622,811,9140,4570,2285,9815,12554,
                   6277,11875,13584,6792,3396,1698,849,9097,13285,15315,16328,8164,4082,2041,8669,
                   13007,15174,7587,11504,5752,2876,1438,719,9030,4515,10992,5496,2748,1374,687,
                   9078,4539,11004,5502,2751,10110,5055,11262,5631,10462,5231,10262,5131,10276,5138,
                   2569,10021,12723,15096,7548,3774,1887,8590,4295,10818,5409,10417,13945,14621,16047,
                   15734,7867,11644,5822,2911,10126,5063,11202,5601,10449,13897,14597,16035,15728,7864,
                   3932,1966,983,9162,4581,10963,14152,7076,3538,1769,8533,12939,15204,7602,3801,
                   9549,12423,14946,7473,11449,13437,14367,15918,7959,11690,5845,10571,13956,6978,3489,
                   9457,12377,14861,16167,15794,7897,11597,13447,14434,7217,11321,13373,14399,15934,7967,
                   11694,5847,10570,5285,10355,13848,6924,3462,1731,8512,4256,2128,1064,532,266,
                   133,8803,13072,6536,3268,1634,817,9145,13309,15327,16334,8167,11730,5865,10581,
                   13963,14692,7346,3673,9485,12455,14962,7481,11453,13439,14366,7183,11302,5651,10536,
                   5268,2634,1317,8371,12920,6460,3230,1615,8454,4227,10848,5424,2712,1356,678,
                   339,8840,4420,2210,1105,8201,12837,15155,16312,8156,4078,2039,8666,4333,10839,
                   14090,7045,12259,13776,6888,3444,1722,861,9103,13286,6643,11992,5996,2998,1499,
                   8396,4198,2099,9784,4892,2446,1223,8258,4129,10801,14137,14781,16127,15710,7855,
                   11638,5819,10620,5310,2655,9998,4999,11234,5617,10457,13901,14599,16034,8017,11657,
                   13541,14419,15880,7940,3970,1985,8641,12993,15169,16257,15841,15569,15433,15365,15395,
                   15408,7704,3852,1926,963,9152,4576,2288,1144,572,286,143,8806,4403,10936,
                   5468,2734,1367,8330,4165,10755,14112,7056,3528,1764,882,441,8957,13151,15246,
                   7623,11458,5729,10513,13993,14709,16027,15724,7862,3931,9612,4806,2403,9872,4936,
                   2468,1234,617,8981,13227,15348,7674,3837,9567,12430,6215,11778,5889,10657,14065,
                   14681,16013,15719,15506,7753,11525,13475,14448,7224,3612,1806,903,9186,4593,10969,
                   14157,14727,16098,8049,11673,13549,14423,15882,7941,11683,13552,6776,3388,1694,847,
                   9094,4547,10944,5472,2736,1368,684,342,171,8820,4410,2205,9839,12566,6283,
                   11876,5938,2969,10221,12759,15050,7525,11411,13416,6708,3354,1677,8551,12946,6473,
                   11909,13667,14480,7240,3620,1810,905,9189,13267,15304,7652,3826,1913,8605,13039,
                   15190,7595,11508,5754,2877,10175,12798,6399,11870,5935,10678,5339,10316,5158,2579,
                   10024,5012,2506,1253,8275,12808,6404,3202,1601,8449,12961,15217,16281,15853,15575,
                   15434,7717,11571,13496,6748,3374,1687,8554,4277,10875,14108,7054,3527,9410,4705,
                   11025,14249,14837,16091,15692,7846,3923,9608,4804,2402,1201,8313,12829,15151,16310,
                   8155,11724,5862,2931,10136,5068,2534,1267,8280,4140,2070,1035,8228,4114,2057,
                   9765,12595,15032,7516,3758,1879,8586,4293,10819,14080,7040,3520,1760,880,440,
                   220,110,55,8762,4381,10927,14198,7099,12284,6142,3071,10206,5103,11222,5611,
                   10452,5226,2613,10043,12732,6366,3183,9238,4619,11044,5522,2761,10053,12675,15072,
                   7536,3768,1884,942,471,8906,4453,10899,14184,7092,3546,1773,8535,12938,6469,
                   11907,13664,6832,3416,1708,854,427,8948,4474,2237,9855,12574,6287,11878,5939,
                   10680,5340,2670,1335,8378,4189,10767,14118,7059,12264,6132,3066,1533,8415,12878,
                   6439,11954,5977,10637,14055,14674,7337,11381,13339,14380,7190,3595,9508,4754,2377,
                   9861,12643,14992,7496,3748,1874,937,9205,13275,15308,7654,3827,9560,4780,2390,
                   1195,8308,4154,2077,9775,12598,6299,11884,5942,2971,10220,5110,2555,9948,4974,
                   2487,9978,4989,11167,14318,7159,12250,6125,10711,14026,7013,12179,13800,6900,3450,
                   1725,8575,12958,6479,11910,5955,10624,5312,2656,1328,664,332,166,83,8712,
                   4356,2178,1089,8193,12833,15153,16313,15869,15583,15438,7719,11570,5785,10605,13975,
                   14698,7349,11387,13340,6670,3335,9378,4689,11017,14245,14835,16088,8044,4022,2011,
                   8652,4326,2163,9752,4876,2438,1219,8256,4128,2064,1032,516,258,129,8801,
                   13073,15273,16373,15835,15564,7782,3891,9656,4828,2414,1207,8314,4157,10815,14142,
                   7071,12270,6135,10714,5357,10327,13834,6917,12195,13808,6904,3452,1726,863,9102,
                   4551,10946,5473,10385,13929,14613,16043,15732,7866,3933,9615,12518,6259,11800,5900,
                   2950,1475,8384,4192,2096,1048,524,262,131,8800,4400,2200,1100,550,275,
                   8872,4436,2218,1109,8203,12836,6418,3209,9317,12307,14888,7444,3722,1861,8579,
                   13024,6512,3256,1628,814,407,8938,4469,10907,14188,7094,3547,9420,4710,2355,
                   9912,4956,2478,1239,8266,4133,10803,14136,7068,3534,1767,8530,4265,10869,14107,
                   14764,7382,3691,9492,4746,2373,9859,12640,6320,3160,1580,790,395,8932,4466,
                   2233,9853,12575,15022,7511,11402,5701,10499,13984,6992,3496,1748,874,437,8955,
                   13148,6574,3287,9290,4645,11059,14264,7132,3566,1783,8538,4269,10871,14106,7053,
                   12263,13778,6889,12117,13707,14564,7282,3641,9533,12479,14974,7487,11454,5727,10510,
                   5255,10338,5169,10297,13885,14655,16062,8031,11662,5831,10562,5281,10353,13849,14637,
                   16055,15738,7869,11647,13470,6735,12038,6019,10720,5360,2680,1340,670,335,8838,
                   4419,10880,5440,2720,1360,680,340,170,85,8715,13092,6546,3273,9285,12291,
                   14880,7440,3720,1860,930,465,8905,13125,15235,16352,8176,4088,2044,1022,511,
                   8926,4463,10902,5451,10372,5186,2593,10033,12729,15101,16223,15758,7879,11586,5793,
                   10609,13977,14701,16023,15722,7861,11643,13468,6734,3367,9394,4697,11021,14247,14834,
                   7417,11357,13327,14374,7187,11304,5652,2826,1413,8419,12880,6440,3220,1610,805,
                   9139,13304,6652,3326,1663,8478,4239,10854,5427,10424,5212,2606,1303,8362,4181,
                   10763,14116,7058,3529,9413,12355,14848,7424,3712,1856,928,464,232,116,58,
                   29,8751,13110,6555,12012,6006,3003,10236,5118,2559,9950,4975,11158,5579,10436,
                   5218,2609,10041,12733,15103,16222,8111,11766,5883,10588,5294,2647,9994,4997,11235,
                   14288,7144,3572,1786,893,9119,13294,6647,11994,5997,10647,14058,7029,12187,13804,
                   6902,3451,9372,4686,2343,9906,4953,11149,14311,14802,7401,11349,13323,14372,7186,
                   3593,9509,12467,14968,7484,3742,1871,8582,4291,10816,5408,2704,1352,676,338,
                   169,8821,13083,15276,7638,3819,9556,4778,2389,9867,12644,6322,3161,9229,12327,
                   14898,7449,11437,13431,14362,7181,11303,13362,6681,12077,13751,14586,7293,11295,13358,
                   6679,12074,6037,10731,14036,7018,3509,9467,12380,6190,3095,9258,4629,11051,14260,
                   7130,3565,9431,12362,6181,11827,13624,6812,3406,1703,8562,4281,10877,14111,14766,
                   7383,11338,5669,10547,14008,7004,3502,1751,8522,4261,10867,14104,7052,3526,1763,
                   8528,4264,2132,1066,533,9003,13236,6618,3309,9303,12298,6149,11811,13616,6808,
                   3404,1702,851,9096,4548,2274,1137,8217,12845,15159,16314,8157,11727,13510,6755,
                   12048,6024,3012,1506,753,9049,13197,15335,16338,8169,11733,13515,14404,7202,3601,
                   9513,12469,14971,16156,8078,4039,9666,4833,11089,14217,14821,16083,15688,7844,3922,
                   1961,8693,13019,15180,7590,3795,9544,4772,2386,1193,8309,12827,15148,7574,3787,
                   9540,4770,2385,9865,12645,14995,16232,8116,4058,2029,8663,13002,6501,11923,13672,
                   6836,3418,1709,8567,12954,6477,11911,13666,6833,12153,13725,14575,15958,7979,11700,
                   5850,2925,10135,12778,6389,11867,13580,6790,3395,9344,4672,2336,1168,584,292,
                   146,73,8709,13091,15280,7640,3820,1910,955,9212,4606,2303,9822,4911,11190,
                   5595,10444,5222,2611,10040,5020,2510,1255,8274,4137,10805,14139,14780,7390,3695,
                   9494,4747,11108,5554,2777,10061,12679,15074,7537,11417,13421,14359,15914,7957,11691,
                   13556,6778,3389,9407,12414,6207,11838,5919,10670,5335,10314,5157,10291,13880,6940,
                   3470,1735,8514,4257,10865,14105,14765,16119,15706,7853,11639,13466,6733,12039,13730,
                   6865,12105,13701,14563,15952,7976,3988,1994,997,9171,13256,6628,3314,1657,8477,
                   12975,15222,7611,11516,5758,2879,10174,5087,11214,5607,10450,5225,10261,13867,14644,
                   7322,3661,9479,12450,6225,11785,13605,14515,15992,7996,3998,1999,8646,4323,10832,
                   5416,2708,1354,677,9075,13208,6604,3302,1651,8472,4236,2118,1059,8240,4120,
                   2060,1030,515,8992,4496,2248,1124,562,281,8877,13175,15258,7629,11463,13378,
                   6689,12081,13753,14589,15967,15630,7815,11618,5809,10617,13981,14703,16022,8011,11652,
                   5826,2913,10129,12777,15061,16203,15748,7874,3937,9617,12521,14933,16139,15780,7890,
                   3945,9621,12523,14932,7466,3733,9579,12436,6218,3109,9267,12344,6172,3086,1543,
                   8482,4241,10857,14101,14763,16116,8058,4029,9727,12510,6255,11798,5899,10660,5330,
                   2665,10005,12715,15092,7546,3773,9599,12446,6223,11782,5891,10656,5328,2664,1332,
                   666,333,8839,13154,6577,12025,13661,14479,15974,7987,11704,5852,2926,1463,8442,
                   4221,10783,14126,7063,12266,6133,10715,14028,7014,3507,9464,4732,2366,1183,8302,
                   4151,10810,5405,10415,13942,6971,12220,6110,3055,10198,5099,11220,5610,2805,10075,
                   12684,6342,3171,9232,4616,2308,1154,577,8961,13217,15345,16345,15821,15559,15426,
                   7713,11569,13497,14461,15903,15662,7831,11626,5813,10619,13980,6990,3495,9458,4729,
                   11037,14255,14838,7419,11356,5678,2839,10154,5077,11211,14276,7138,3569,9433,12365,
                   14855,16162,8081,11753,13525,14411,15876,7938,3969,9697,12497,14921,16133,15779,15600,
                   7800,3900,1950,975,9158,4579,10960,5480,2740,1370,685,9079,13210,6605,11975,
                   13634,6817,12145,13721,14573,15959,15626,7813,11619,13456,6728,3364,1682,841,9093,
                   13283,15312,7656,3828,1914,957,9215,13278,6639,11990,5995,10644,5322,2661,10003,
                   12712,6356,3178,1589,8507,12988,6494,3247,9334,4667,11068,5534,2767,10054,5027,
                   11248,5624,2812,1406,703,9086,4543,11006,5503,10398,5199,10246,5123,10272,5136,
                   2568,1284,642,321,8833,13153,15249,16361,15829,15563,15428,7714,3857,9641,12533,
                   14939,16140,8070,4035,9664,4832,2416,1208,604,302,151,8810,4405,10939,14204,
                   7102,3551,9422,4711,11026,5513,10469,13907,14600,7300,3650,1825,8625,13049,15197,
                   16271,15846,7923,11608,5804,2902,1451,8436,4218,2109,9791,12606,6303,11886,5943,
                   10682,5341,10319,13830,6915,12192,6096,3048,1524,762,381,8863,13166,6583,12026,
                   6013,10655,14062,7031,12186,6093,10695,14018,7009,12177,13801,14549,15947,15620,7810,
                   3905,9601,12513,14929,16137,15781,15603,15448,7724,3862,1931,8676,4338,2169,9757,
                   12591,15030,7515,11404,5702,2851,10160,5080,2540,1270,635,8988,4494,2247,9794,
                   4897,11185,14329,14813,16079,15686,7843,11632,5816,2908,1454,727,9034,4517,10995,
                   14168,7084,3542,1771,8532,4266,2133,9739,12580,6290,3145,9221,12323,14896,7448,
                   3724,1862,931,9200,4600,2300,1150,575,9022,4511,10990,5495,10394,5197,10247,
                   13858,6929,12201,13813,14555,15948,7974,3987,9704,4852,2426,1213,8319,12830,6415,
                   11942,5971,10632,5316,2658,1329,8377,12925,15135,16302,8151,11722,5861,10579,13960,
                   6980,3490,1745,8521,12933,15203,16272,8136,4068,2034,1017,9181,13263,15302,7651,
                   11472,5736,2868,1434,717,9031,13186,6593,11969,13633,14465,15969,15633,15529,15477,
                   15387,15404,7702,3851,9636,4818,2409,9877,12651,14996,7498,3749,9587,12440,6220,
                   3110,1555,8488,4244,2122,1061,8243,12856,6428,3214,1607,8450,4225,10849,14097,
                   14761,16117,15707,15500,7750,3875,9648,4824,2412,1206,603,8972,4486,2243,9792,
                   4896,2448,1224,612,306,153,8813,13079,15274,7637,11467,13380,6690,3345,9385,
                   12405,14875,16172,8086,4043,9668,4834,2417,9881,12653,14999,16234,8117,11771,13532,
                   6766,3383,9402,4701,11023,14246,7123,12232,6116,3058,1529,8413,12879,15110,7555,
                   11488,5744,2872,1436,718,359,8850,4425,10885,14179,14736,7368,3684,1842,921,
                   9197,13271,15306,7653,11475,13384,6692,3346,1673,8549,12947,15208,7604,3802,1901,
                   8599,13034,6517,11931,13676,6838,3419,9356,4678,2339,9904,4952,2476,1238,619,
                   8980,4490,2245,9795,12544,6272,3136,1568,784,392,196,98,49,8761,13117,
                   15295,16382,8191,11742,5871,10582,5291,10356,5178,2589,10031,12726,6363,11852,5926,
                   2963,10216,5108,2554,1277,8287,12814,6407,11938,5969,10633,14053,14675,16008,8004,
                   4002,2001,8649,12997,15171,16256,8128,4064,2032,1016,508,254,127,8734,4367,
                   10918,5459,10376,5188,2594,1297,8361,12917,15131,16300,8150,4075,9684,4842,2421,
                   9883,12652,6326,3163,9228,4614,2307,9888,4944,2472,1236,618,309,8891,13180,
                   6590,3295,9294,4647,11058,5529,10477,13911,14602,7301,11363,13328,6664,3332,1666,
                   833,9089,13281,15313,16329,15813,15555,15424,7712,3856,1928,964,482,241,8793,
                   13069,15271,16370,8185,11741,13519,14406,7203,11312,5656,2828,1414,707,9024,4512,
                   2256,1128,564,282,141,8807,13074,6537,12005,13651,14472,7236,3618,1809,8617,
                   13045,15195,16268,8134,4067,9680,4840,2420,1210,605,8975,13222,6611,11976,5988,
                   2994,1497,8397,12871,15106,7553,11489,13393,14345,15909,15667,15544,7772,3886,1943,
                   8682,4341,10843,14092,7046,3523,9408,4704,2352,1176,588,294,147,8808,4404,
                   2202,1101,8199,12834,6417,11945,13685,14491,15980,7990,3995,9708,4854,2427,9884,
                   4942,2471,9970,4985,11165,14319,14806,7403,11348,5674,2837,10155,12788,6394,3197,
                   9247,12334,6167,11818,5909,10667,14068,7034,3517,9471,12382,6191,11830,5915,10668,
                   5334,2667,10004,5002,2501,9923,12608,6304,3152,1576,788,394,197,8771,13056,
                   6528,3264,1632,816,408,204,102,51,8760,4380,2190,1095,8194,4097,10785,
                   14129,14777,16125,15711,15502,7751,11522,5761,10593,13969,14697,16021,15723,15508,7754,
                   3877,9651,12536,6268,3134,1567,8494,4247,10858,5429,10427,13948,6974,3487,9454,
                   4727,11034,5517,10471,13906,6953,12213,13819,14556,7278,3639,9530,4765,11119,14230,
                   7115,12228,6114,3057,10201,12749,15047,16194,8097,11761,13529,14413,15879,15650,7825,
                   11625,13461,14443,15892,7946,3973,9699,12496,6248,3124,1562,781,9127,13298,6649,
                   11997,13647,14470,7235,11264,5632,2816,1408,704,352,176,88,44,22,11,
                   8740,4370,2185,9829,12563,15016,7508,3754,1877,8587,13028,6514,3257,9341,12319,
                   14894,7447,11434,5717,10507,13988,6994,3497,9461,12379,14860,7430,3715,9568,4784,
                   2392,1196,598,299,8884,4442,2221,9847,12570,6285,11879,13586,6793,12133,13715,
                   14568,7284,3642,1821,8623,13046,6523,11932,5966,2983,10226,5113,11229,14287,14790,
                   7395,11344,5672,2836,1418,709,9027,13184,6592,3296,1648,824,412,206,103,
                   8722,4361,10917,14195,14744,7372,3686,1843,8632,4316,2158,1079,8250,4125,10799,
                   14134,7067,12268,6134,3067,10204,5102,2551,9946,4973,11159,14314,7157,12251,13772,
                   6886,3443,9368,4684,2342,1171,8296,4148,2074,1037,8231,12850,6425,11949,13687,
                   14490,7245,11271,13346,6673,12073,13749,14587,15964,7982,3991,9706,4853,11099,14220,
                   7110,3555,9424,4712,2356,1178,589,8967,13218,6609,11977,13637,14467,15968,7984,
                   3992,1996,998,499,8920,4460,2230,1115,8204,4102,2051,9760,4880,2440,1220,
                   610,305,8889,13181,15263,16366,8183,11738,5869,10583,13962,6981,12163,13792,6896,
                   3448,1724,862,431,8950,4475,10908,5454,2727,10098,5049,11261,14303,14798,7399,
                   11346,5673,10549,14011,14716,7358,3679,9486,4743,11106,5553,10489,13917,14607,16038,
                   8019,11656,5828,2914,1457,8441,12893,15119,16294,8147,11720,5860,2930,1465,8445,
                   12895,15118,7559,11490,5745,10521,13997,14711,16026,8013,11655,13538,6769,12057,13741,
                   14583,15962,7981,11703,13562,6781,12063,13742,6871,12106,6053,10739,14040,7020,3510,
                   1755,8524,4262,2131,9736,4868,2434,1217,8257,12801,15137,16305,15865,15581,15439,
                   15366,7683,11552,5776,2888,1444,722,361,8853,13163,15252,7626,3813,9555,12424,
                   6212,3106,1553,8489,12981,15227,16284,8142,4071,9682,4841,11093,14219,14820,7410,
                   3705,9501,12463,14966,7483,11452,5726,2863,10166,5083,11212,5606,2803,10072,5036,
                   2518,1259,8276,4138,2069,9771,12596,6298,3149,9223,12322,6161,11817,13621,14523,
                   15996,7998,3999,9710,4855,11098,5549,10487,13914,6957,12215,13818,6909,12127,13710,
                   6855,12098,6049,10737,14041,14669,16007,15714,7857,11641,13469,14447,15894,7947,11684,
                   5842,2921,10133,12779,15060,7530,3765,9595,12444,6222,3111,9266,4633,11053,14263,
                   14842,7421,11359,13326,6663,12066,6033,10729,14037,14667,16004,8002,4001,9713,12505,
                   14925,16135,15778,7889,11593,13445,14435,15888,7944,3972,1986,993,9169,13257,15301,
                   16323,15808,7904,3952,1976,988,494,247,8794,4397,10935,14202,7101,12287,13790,
                   6895,12118,6059,10740,5370,2685,10015,12718,6359,11850,5925,10675,14072,7036,3518,
                   1759,8526,4263,10866,5433,10429,13951,14622,7311,11366,5683,10552,5276,2638,1319,
                   8370,4185,10765,14119,14770,7385,11341,13319,14370,7185,11305,13365,14395,15932,7966,
                   3983,9702,4851,11096,5548,2774,1387,8340,4170,2085,9779,12600,6300,3150,1575,
                   8498,4249,10861,14103,14762,7381,11339,13316,6658,3329,9377,12401,14873,16173,15799,
                   15610,7805,11551,13486,6743,12042,6021,10723,14032,7016,3508,1754,877,9111,13290,
                   6645,11995,13644,6822,3411,9352,4676,2338,1169,8297,12821,15147,16308,8154,4077,
                   9687,12490,6245,11795,13608,6804,3402,1701,8563,12952,6476,3238,1619,8456,4228,
                   2114,1057,8241,12857,15165,16319,15870,7935,11614,5807,10614,5307,10364,5182,2591,
                   10030,5015,11242,5621,10459,13900,6950,3475,9448,4724,2362,1181,8303,12822,6411,
                   11940,5970,2985,10229,12763,15052,7526,3763,9592,4796,2398,1199,8310,4155,10812,
                   5406,2703,10086,5043,11256,5628,2814,1407,8350,4175,10758,5379,10400,5200,2600,
                   1300,650,325,8835,13152,6576,3288,1644,822,411,8940,4470,2235,9852,4926,
                   2463,9966,4983,11162,5581,10439,13890,6945,12209,13817,14557,15951,15622,7811,11616,
                   5808,2904,1452,726,363,8852,4426,2213,9843,12568,6284,3142,1571,8496,4248,
                   2124,1062,531,9000,4500,2250,1125,8211,12840,6420,3210,1605,8451,12960,6480,
                   3240,1620,810,405,8939,13140,6570,3285,9291,12292,6146,3073,9249,12337,14905,
                   16189,15807,15614,7807,11550,5775,10598,5299,10360,5180,2590,1295,8358,4179,10760,
                   5380,2690,1345,8321,12897,15121,16297,15861,15579,15436,7718,3859,9640,4820,2410,
                   1205,8315,12828,6414,3207,9314,4657,11065,14269,14847,16094,8047,11670,5835,10564,
                   5282,2641,9993,12709,15091,16216,8108,4054,2027,8660,4330,2165,9755,12588,6294,
                   3147,9220,4610,2305,9889,12657,15001,16237,15767,15594,7797,11547,13484,6742,3371,
                   9396,4698,2349,9911,12666,6333,11903,13598,6799,12134,6067,10744,5372,2686,1343,
                   8382,4191,10766,5383,10402,5201,10249,13861,14643,16056,8028,4014,2007,8650,4325,
                   10835,14088,7044,3522,1761,8529,12937,15205,16275,15848,7924,3962,1981,8703,13022,
                   6511,11926,5963,10628,5314,2657,10001,12713,15093,16219,15756,7878,3939,9616,4808,
                   2404,1202,601,8973,13223,15346,7673,11485,13391,14342,7171,11296,5648,2824,1412,
                   706,353,8849,13161,15253,16363,15828,7914,3957,9627,12524,6262,3131,9276,4638,
                   2319,9894,4947,11144,5572,2786,1393,8345,12909,15127,16298,8149,11723,13508,6754,
                   3377,9401,12413,14879,16174,8087,11754,5877,10587,13964,6982,3491,9456,4728,2364,
                   1182,591,8966,4483,10976,5488,2744,1372,686,343,8842,4421,10883,14176,7088,
                   3544,1772,886,443,8956,4478,2239,9854,4927,11198,5599,10446,5223,10258,5129,
                   10277,13875,14648,7324,3662,1831,8626,4313,10829,14087,14754,7377,11337,13317,14371,
                   15920,7960,3980,1990,995,9168,4584,2292,1146,573,9023,13246,6623,11982,5991,
                   10642,5321,10309,13827,14624,7312,3656,1828,914,457,8901,13123,15232,7616,3808,
                   1904,952,476,238,119,8730,4365,10919,14194,7097,12285,13791,14542,7271,11282,
                   5641,10533,14003,14712,7356,3678,1839,8630,4315,10828,5414,2707,10088,5044,2522,
                   1261,8279,12810,6405,11939,13680,6840,3420,1710,855,9098,4549,10947,14144,7072,
                   3536,1768,884,442,221,8783,13062,6531,12000,6000,3000,1500,750,375,8858,
                   4429,10887,14178,7089,12281,13789,14543,15942,7971,11696,5848,2924,1462,731,9036,
                   4518,2259,9800,4900,2450,1225,8261,12803,15136,7568,3784,1892,946,473,8909,
                   13127,15234,7617,11457,13377,14337,15905,15665,15545,15485,15391,15406,7703,11562,5781,
                   10603,13972,6986,3493,9459,12376,6188,3094,1547,8484,4242,2121,9733,12579,15024,
                   7512,3756,1878,939,9204,4602,2301,9823,12558,6279,11874,5937,10681,14077,14687,
                   16014,8007,11650,5825,10561,13953,14689,16017,15721,15509,15467,15380,7690,3845,9635,
                   12528,6264,3132,1566,783,9126,4563,10952,5476,2738,1369,8333,12903,15122,7561,
                   11493,13395,14344,7172,3586,1793,8609,13041,15193,16269,15847,15570,7785,11541,13483,
                   14452,7226,3613,9519,12470,6235,11788,5894,2947,10208,5104,2552,1276,638,319,
                   8894,4447,10894,5447,10370,5185,10241,13857,14641,16057,15741,15519,15470,7735,11578,
                   5789,10607,13974,6987,12164,6082,3041,10193,12745,15045,16195,15744,7872,3936,1968,
                   984,492,246,123,8732,4366,2183,9826,4913,11193,14333,14815,16078,8039,11666,
                   5833,10565,13955,14688,7344,3672,1836,918,459,8900,4450,2225,9849,12573,15023,
                   16246,8123,11772,5886,2943,10142,5071,11206,5603,10448,5224,2612,1306,653,9063,
                   13202,6601,11973,13635,14464,7232,3616,1808,904,452,226,113,8729,13101,15287,
                   16378,8189,11743,13518,6759,12050,6025,10725,14035,14664,7332,3666,1833,8629,13051,
                   15196,7598,3799,9546,4773,11123,14232,7116,3558,1779,8536,4268,2134,1067,8244,
                   4122,2061,9767,12594,6297,11885,13591,14506,7253,11275,13348,6674,3337,9381,12403,
                   14872,7436,3718,1859,8576,4288,2144,1072,536,268,134,67,8704,4352,2176,
                   1088,544,272,136,68,34,17,8745,13109,15291,16380,8190,4095,9694,4847,
                   11094,5547,10484,5242,2621,10047,12734,6367,11854,5927,10674,5337,10317,13831,14626,
                   7313,11369,13333,14379,15924,7962,3981,9703,12498,6249,11797,13611,14516,7258,3629,
                   9527,12474,6237,11791,13606,6803,12136,6068,3034,1517,8407,12874,6437,11955,13688,
                   6844,3422,1711,8566,4283,10876,5438,2719,10094,5047,11258,5629,10463,13902,6951,
                   12210,6105,10701,14023,14658,7329,11377,13337,14381,15927,15674,7837,11631,13462,6731,
                   12036,6018,3009,10177,12737,15041,16193,15745,15585,15441,15369,15397,15411,15416,7708,
                   3854,1927,8674,4337,10841,14093,14759,16114,8057,11677,13551,14422,7211,11316,5658,
                   2829,10151,12786,6393,11869,13583,14502,7251,11272,5636,2818,1409,8417,12881,15113,
                   16293,15859,15576,7788,3894,1947,8684,4342,2171,9756,4878,2439,9954,4977,11161,
                   14317,14807,16074,8037,11667,13544,6772,3386,1693,8559,12950,6475,11908,5954,2977,
                   10225,12761,15053,16199,15746,7873,11585,13441,14433,15889,15657,15541,15483,15388,7694,
                   3847,9634,4817,11081,14213,14819,16080,8040,4020,2010,1005,9175,13258,6629,11987,
                   13640,6820,3410,1705,8565,12955,15212,7606,3803,9548,4774,2387,9864,4932,2466,
                   1233,8265,12805,15139,16304,8152,4076,2038,1019,9180,4590,2295,9818,4909,11191,
                   14330,7165,12255,13774,6887,12114,6057,10741,14043,14668,7334,3667,9480,4740,2370,
                   1185,8305,12825,15149,16311,15866,7933,11615,13454,6727,12034,6017,10721,14033,14665,
                   16005,15715,15504,7752,3876,1938,969,9157,13251,15296,7648,3824,1912,956,478,
                   239,8790,4395,10932,5466,2733,10103,12698,6349,11847,13570,6785,12129,13713,14569,
                   15957,15627,15524,7762,3881,9653,12539,14940,7470,3735,9578,4789,11131,14236,7118,
                   3559,9426,4713,11029,14251,14836,7418,3709,9503,12462,6231,11786,5893,10659,14064,
                   7032,3516,1758,879,9110,4555,10948,5474,2737,10105,12701,15087,16214,8107,11764,
                   5882,2941,10143,12782,6391,11866,5933,10679,14074,7037,12191,13806,6903,12122,6061,
                   10743,14042,7021,12183,13802,6901,12123,13708,6854,3427,9360,4680,2340,1170,585,
                   8965,13219,15344,7672,3836,1918,959,9214,4607,10974,5487,10390,5195,10244,5122,
                   2561,10017,12721,15097,16221,15759,15590,7795,11544,5772,2886,1443,8432,4216,2108,
                   1054,527,8998,4499,10984,5492,2746,1373,8335,12902,6451,11960,5980,2990,1495,
                   8394,4197,10771,14120,7060,3530,1765,8531,12936,6468,3234,1617,8457,12965,15219,
                   16280,8140,4070,2035,8664,4332,2166,1083,8252,4126,2063,9766,4883,11176,5588,
                   2794,1397,8347,12908,6454,3227,9324,4662,2331,9900,4950,2475,9972,4986,2493,
                   9983,12638,6319,11894,5947,10684,5342,2671,10006,5003,11236,5618,2809,10077,12687,
                   15078,7539,11416,5708,2854,1427,8424,4212,2106,1053,8239,12854,6427,11948,5974,
                   2987,10228,5114,2557,9951,12622,6311,11890,5945,10685,14079,14686,7343,11382,5691,
                   10556,5278,2639,9990,4995,11232,5616,2808,1404,702,351,8846,4423,10882,5441,
                   10369,13921,14609,16041,15733,15515,15468,7734,3867,9644,4822,2411,9876,4938,2469,
                   9971,12632,6316,3158,1579,8500,4250,2125,9735,12578,6289,11881,13589,14507,15988,
                   7994,3997,9711,12502,6251,11796,5898,2949,10211,12752,6376,3188,1594,797,9135,
                   13302,6651,11996,5998,2999,10234,5117,11231,14286,7143,12242,6121,10709,14027,14660,
                   7330,3665,9481,12453,14963,16152,8076,4038,2019,8656,4328,2164,1082,541,9007,
                   13238,6619,11980,5990,2995,10232,5116,2558,1279,8286,4143,10806,5403,10412,5206,
                   2603,10036,5018,2509,9927,12610,6305,11889,13593,14509,15991,15642,7821,11623,13458,
                   6729,12037,13731,14576,7288,3644,1822,911,9190,4595,10968,5484,2742,1371,8332,
                   4166,2083,9776,4888,2444,1222,611,8976,4488,2244,1122,561,9017,13245,15359,
                   16350,8175,11734,5867,10580,5290,2645,9995,12708,6354,3177,9237,12331,14900,7450,
                   3725,9575,12434,6217,11781,13603,14512,7256,3628,1814,907,9188,4594,2297,9821,
                   12559,15014,7507,11400,5700,2850,1425,8425,12885,15115,16292,8146,4073,9685,12491,
                   14916,7458,3729,9577,12437,14955,16148,8074,4037,9667,12480,6240,3120,1560,780,
                   390,195,8768,4384,2192,1096,548,274,137,8805,13075,15272,7636,3818,1909,
                   8603,13036,6518,3259,9340,4670,2335,9902,4951,11146,5573,10435,13888,6944,3472,
                   1736,868,434,217,8781,13063,15266,7633,11465,13381,14339,15904,7952,3976,1988,
                   994,497,8921,13133,15239,16354,8177,11737,13517,14407,15874,7937,11681,13553,14425,
                   15885,15655,15538,7769,11533,13479,14450,7225,11325,13375,14398,7199,11310,5655,10538,
                   5269,10347,13844,6922,3461,9443,12368,6184,3092,1546,773,9123,13296,6648,3324,
                   1662,831,9150,4575,10958,5479,10386,5193,10245,13859,14640,7320,3660,1830,915,
                   9192,4596,2298,1149,8223,12846,6423,11946,5973,10635,14052,7026,3513,9469,12383,
                   14862,7431,11426,5713,10505,13989,14707,16024,8012,4006,2003,8648,4324,2162,1081,
                   8253,12863,15166,7583,11502,5751,10522,5261,10343,13842,6921,12197,13811,14552,7276,
                   3638,1819,8620,4310,2155,9748,4874,2437,9955,12624,6312,3156,1578,789,9131,
                   13300,6650,3325,9311,12302,6151,11810,5905,10665,14069,14683,16012,8006,4003,9712,
                   4856,2428,1214,607,8974,4487,10978,5489,10393,13933,14615,16042,8021,11659,13540,
                   6770,3385,9405,12415,14878,7439,11430,5715,10504,5252,2626,1313,8369,12921,15133,
                   16303,15862,7931,11612,5806,2903,10122,5061,11203,14272,7136,3568,1784,892,446,
                   223,8782,4391,10930,5465,10381,13927,14610,7305,11365,13331,14376,7188,3594,1797,
                   8611,13040,6520,3260,1630,815,9142,4571,10956,5478,2739,10104,5052,2526,1263,
                   8278,4139,10804,5402,2701,10087,12690,6345,11845,13571,14496,7248,3624,1812,906,
                   453,8899,13120,6560,3280,1640,820,410,205,8775,13058,6529,12001,13649,14473,
                   15973,15635,15528,7764,3882,1941,8683,13012,6506,3253,9339,12316,6158,3079,9250,
                   4625,11049,14261,14843,16092,8046,4023,9722,4861,11103,14222,7111,12226,6113,10705,
                   14025,14661,16003,15712,7856,3928,1964,982,491,8916,4458,2229,9851,12572,6286,
                   3143,9218,4609,11041,14257,14841,16093,15695,15494,7747,11520,5760,2880,1440,720,
                   360,180,90,45,8759,13114,6557,12015,13654,6827,12148,6074,3037,10191,12742,
                   6371,11856,5928,2964,1482,741,9043,13192,6596,3298,1649,8473,12973,15223,16282,
                   8141,11719,13506,6753,12049,13737,14581,15963,15628,7814,3907,9600,4800,2400,1200,
                   600,300,150,75,8708,4354,2177,9825,12561,15017,16245,15771,15596,7798,3899,
                   9660,4830,2415,9878,4939,11140,5570,2785,10065,12681,15077,16211,15752,7876,3938,
                   1969,8697,13021,15183,16262,8131,11712,5856,2928,1464,732,366,183,8826,4413,
                   10943,14206,7103,12286,6143,10718,5359,10326,5163,10292,5146,2573,10023,12722,6361,
                   11853,13575,14498,7249,11273,13349,14387,15928,7964,3982,1991,8642,4321,10833,14089,
                   14757,16115,15704,7852,3926,1963,8692,4346,2173,9759,12590,6295,11882,5941,10683,
                   14076,7038,3519,9470,4735,11038,5519,10470,5235,10264,5132,2566,1283,8352,4176,
                   2088,1044,522,261,8867,13168,6584,3292,1646,823,9146,4573,10959,14150,7075,
                   12272,6136,3068,1534,767,9054,4527,10998,5499,10396,5198,2599,10034,5017,11245,
                   14295,14794,7397,11347,13320,6660,3330,1665,8545,12945,15209,16277,15851,15572,7786,
                   3893,9659,12540,6270,3135,9278,4639,11054,5527,10474,5237,10267,13868,6934,3467,
                   9444,4722,2361,9917,12671,15006,7503,11398,5699,10496,5248,2624,1312,656,328,
                   164,82,41,8757,13115,15292,7646,3823,9558,4779,11124,5562,2781,10063,12678,
                   6339,11840,5920,2960,1480,740,370,185,8829,13087,15278,7639,11466,5733,10515,
                   13992,6996,3498,1749,8523,12932,6466,3233,9329,12313,14893,16183,15802,7901,11599,
                   13446,6723,12032,6016,3008,1504,752,376,188,94,47,8758,4379,10924,5462,
                   2731,10100,5050,2525,9935,12614,6307,11888,5944,2972,1486,743,9042,4521,10997,
                   14171,14732,7366,3683,9488,4744,2372,1186,593,8969,13221,15347,16344,8172,4086,
                   2043,8668,4334,2167,9754,4877,11175,14322,7161,12253,13775,14534,7267,11280,5640,
                   2820,1410,705,9025,13185,15329,16337,15817,15557,15427,15360,7680,3840,1920,960,
                   480,240,120,60,30,15,8742,4371,10920,5460,2730,1365,8331,12900,6450,
                   3225,9325,12311,14890,7445,11435,13428,6714,3357,9391,12406,6203,11836,5918,2959,
                   10214,5107,11224,5612,2806,1403,8348,4174,2087,9778,4889,11181,14327,14810,7405,
                   11351,13322,6661,12067,13744,6872,3436,1718,859,9100,4550,2275,9808,4904,2452,
                   1226,613,8979,13224,6612,3306,1653,8475,12972,6486,3243,9332,4666,2333,9903,
                   12662,6331,11900,5950,2975,10222,5111,11226,5613,10455,13898,6949,12211,13816,6908,
                   3454,1727,8574,4287,10878,5439,10430,5215,10254,5127,10274,5137,10281,13877,14651,
                   16060,8030,4015,9718,4859,11100,5550,2775,10058,5029,11251,14296,7148,3574,1787,
                   8540,4270,2135,9738,4869,11171,14320,7160,3580,1790,895,9118,4559,10950,5475,
                   10384,5192,2596,1298,649,9061,13203,15336,7668,3834,1917,8607,13038,6519,11930,
                   5965,10631,14050,7025,12185,13805,14551,15946,7973,11699,13560,6780,3390,1695,8558,
                   4279,10874,5437,10431,13950,6975,12222,6111,10702,5351,10322,5161,10293,13883,14652,
                   7326,3663,9478,4739,11104,5552,2776,1388,694,347,8844,4422,2211,9840,4920,
                   2460,1230,615,8978,4489,10981,14163,14728,7364,3682,1841,8633,13053,15199,16270,
                   8135,11714,5857,10577,13961,14693,16019,15720,7860,3930,1965,8695,13018,6509,11927,
                   13674,6837,12155,13724,6862,3431,9362,4681,11013,14243,14832,7416,3708,1854,927,
                   9198,4599,10970,5485,10391,13930,6965,12219,13820,6910,3455,9374,4687,11014,5507,
                   10464,5232,2616,1308,654,327,8834,4417,10881,14177,14737,16105,15701,15499,15460,
                   7730,3865,9645,12535,14938,7469,11447,13434,6717,12095,13758,6879,12110,6055,10738,
                   5369,10333,13839,14630,7315,11368,5684,2842,1421,8423,12882,6441,11957,13691,14492,
                   7246,3623,9522,4761,11117,14231,14826,7413,11355,13324,6662,3331,9376,4688,2344,
                   1172,586,293,8883,13176,6588,3294,1647,8470,4235,10852,5426,2713,10093,12695,
                   15082,7541,11419,13420,6710,3355,9388,4694,2347,9908,4954,2477,9975,12634,6317,
                   11895,13594,6797,12135,13714,6857,12101,13699,14560,7280,3640,1820,910,455,8898,
                   4449,10897,14185,14741,16107,15700,7850,3925,9611,12516,6258,3129,9277,12351,14910,
                   7455,11438,5719,10506,5253,10339,13840,6920,3460,1730,865,9105,13289,15317,16331,
                   15812,7906,3953,9625,12525,14935,16138,8069,11747,13520,6760,3380,1690,845,9095,
                   13282,6641,11993,13645,14471,15970,7985,11705,13565,14431,15886,7943,11682,5841,10569,
                   13957,14691,16016,8008,4004,2002,1001,9173,13259,15300,7650,3825,9561,12429,14951,
                   16146,8073,11749,13523,14408,7204,3602,1801,8613,13043,15192,7596,3798,1899,8596,
                   4298,2149,9747,12584,6292,3146,1573,8499,12984,6492,3246,1623,8458,4229,10851,
                   14096,7048,3524,1762,881,9113,13293,15319,16330,8165,11731,13512,6756,3378,1689,
                   8557,12951,15210,7605,11515,13404,6702,3351,9386,4693,11019,14244,7122,3561,9429,
                   12363,14852,7426,3713,9569,12433,14953,16149,15787,15604,7802,3901,9663,12542,6271,
                   11806,5903,10662,5331,10312,5156,2578,1289,8357,12915,15128,7564,3782,1891,8592,
                   4296,2148,1074,537,9005,13239,15354,7677,11487,13390,6695,12082,6041,10733,14039,
                   14666,7333,11379,13336,6668,3334,1667,8544,4272,2136,1068,534,267,8868,4434,
                   2217,9845,12571,15020,7510,3755,9588,4794,2397,9871,12646,6323,11896,5948,2974,
                   1487,8390,4195,10768,5384,2692,1346,673,9073,13209,15341,16343,15818,7909,11603,
                   13448,6724,3362,1681,8553,12949,15211,16276,8138,4069,9683,12488,6244,3122,1561,
                   8493,12983,15226,7613,11519,13406,6703,12086,6043,10732,5366,2683,10012,5006,2503,
                   9922,4961,11153,14313,14805,16075,15684,7842,3921,9609,12517,14931,16136,8068,4034,
                   2017,8657,13001,15173,16259,15840,7920,3960,1980,990,495,8918,4459,10900,5450,
                   2725,10099,12696,6348,3174,1587,8504,4252,2126,1063,8242,4121,10797,14135,14778,
                   7389,11343,13318,6659,12064,6032,3016,1508,754,377,8861,13167,15254,7627,11460,
                   5730,2865,10169,12797,15071,16206,8103,11762,5881,10589,13967,14694,7347,11384,5692,
                   2846,1423,8422,4211,10776,5388,2694,1347,8320,4160,2080,1040,520,260,130,
                   65,8705,13089,15281,16377,15837,15567,15430,7715,11568,5784,2892,1446,723,9032,
                   4516,2258,1129,8213,12843,15156,7578,3789,9543,12418,6209,11777,13601,14513,15993,
                   15645,15535,15478,7739,11580,5790,2895,10118,5059,11200,5600,2800,1400,700,350,
                   175,8822,4411,10940,5470,2735,10102,5051,11260,5630,2815,10078,5039,11254,5627,
                   10460,5230,2615,10042,5021,11247,14294,7147,12244,6122,3061,10203,12748,6374,3187,
                   9240,4620,2310,1155,8288,4144,2072,1036,518,259,8864,4432,2216,1108,554,
                   277,8875,13172,6586,3293,9295,12294,6147,11808,5904,2952,1476,738,369,8857,
                   13165,15255,16362,8181,11739,13516,6758,3379,9400,4700,2350,1175,8298,4149,10811,
                   14140,7070,3535,9414,4707,11024,5512,2756,1378,689,9081,13213,15343,16342,8171,
                   11732,5866,2933,10139,12780,6390,3195,9244,4622,2311,9890,4945,11145,14309,14803,
                   16072,8036,4018,2009,8653,12999,15170,7585,11505,13401,14349,15911,15666,7833,11629,
                   13463,14442,7221,11323,13372,6686,3343,9382,4691,11016,5508,2754,1377,8337,12905,
                   15125,16299,15860,7930,3965,9631,12526,6263,11802,5901,10663,14066,7033,12189,13807,
                   14550,7275,11284,5642,2821,10147,12784,6392,3196,1598,799,9134,4567,10954,5477,
                   10387,13928,6964,3482,1741,8519,12930,6465,11905,13665,14481,15977,15637,15531,15476,
                   7738,3869,9647,12534,6267,11804,5902,2951,10210,5105,11225,14285,14791,16066,8033,
                   11665,13545,14421,15883,15652,7826,3913,9605,12515,14928,7464,3732,1866,933,9203,
                   13272,6636,3318,1659,8476,4238,2119,9730,4865,11169,14321,14809,16077,15687,15490,
                   7745,11521,13473,14449,15897,15661,15543,15482,7741,11583,13502,6751,12046,6023,10722,
                   5361,10329,13837,14631,16050,8025,11661,13543,14418,7209,11317,13371,14396,7198,3599,
                   9510,4755,11112,5556,2778,1389,8343,12906,6453,11963,13692,6846,3423,9358,4679,
                   11010,5505,10465,13905,14601,16037,15731,15512,7756,3878,1939,8680,4340,2170,1085,
                   8255,12862,6431,11950,5975,10634,5317,10307,13824,6912,3456,1728,864,432,216,
                   108,54,27,8748,4374,2187,9828,4914,2457,9965,12631,14986,7493,11395,13408,
                   6704,3352,1676,838,419,8944,4472,2236,1118,559,9014,4507,10988,5494,2747,
                   10108,5054,2527,9934,4967,11154,5577,10437,13891,14592,7296,3648,1824,912,456,
                   228,114,57,8765,13119,15294,7647,11470,5735,10514,5257,10341,13843,14632,7316,
                   3658,1829,8627,13048,6524,3262,1631,8462,4231,10850,5425,10425,13949,14623,16046,
                   8023,11658,5829,10563,13952,6976,3488,1744,872,436,218,109,8727,13098,6549,
                   12011,13652,6826,3413,9355,12388,6194,3097,9261,12343,14906,7453,11439,13430,6715,
                   12092,6046,3023,10182,5091,11216,5608,2804,1402,701,9087,13214,6607,11974,5987,
                   10640,5320,2660,1330,665,9069,13207,15338,7669,11483,13388,6694,3347,9384,4692,
                   2346,1173,8299,12820,6410,3205,9315,12304,6152,3076,1538,769,9121,13297,15321,
                   16333,15815,15554,7777,11537,13481,14453,15899,15660,7830,3915,9604,4802,2401,9873,
                   12649,14997,16235,15764,7882,3941,9619,12520,6260,3130,1565,8495,12982,6491,11916,
                   5958,2979,10224,5112,2556,1278,639,8990,4495,10982,5491,10392,5196,2598,1299,
                   8360,4180,2090,1045,8235,12852,6426,3213,9319,12306,6153,11813,13619,14520,7260,
                   3630,1815,8618,4309,10827,14084,7042,3521,9409,12353,14849,16161,15793,15609,15453,
                   15375,15398,7699,11560,5780,2890,1445,8435,12888,6444,3222,1611,8452,4226,2113,
                   9729,12577,15025,16249,15773,15599,15446,7723,11572,5786,2893,10119,12770,6385,11865,
                   13581,14503,15986,7993,11709,13567,14430,7215,11318,5659,10540,5270,2635,9988,4994,
                   2497,9921,12609,14977,16225,15761,15593,15445,15371,15396,7698,3849,9637,12531,14936,
                   7468,3734,1867,8580,4290,2145,9745,12585,15029,16251,15772,7886,3943,9618,4809,
                   11077,14211,14816,7408,3704,1852,926,463,8902,4451,10896,5448,2724,1362,681,
                   9077,13211,15340,7670,3835,9564,4782,2391,9866,4933,11139,14304,7152,3576,1788,
                   894,447,8958,4479,10910,5455,10374,5187,10240,5120,2560,1280,640,320,160,
                   80,40,20,10,5,8739,13104,6552,3276,1638,819,9144,4572,2286,1143,
                   8218,4109,10791,14130,7065,12269,13783,14538,7269,11283,13352,6676,3338,1669,8547,
                   12944,6472,3236,1618,809,9141,13307,15324,7662,3831,9562,4781,11127,14234,7117,
                   12231,13762,6881,12113,13705,14565,15955,15624,7812,3906,1953,8689,13017,15181,16263,
                   15842,7921,11609,13453,14439,15890,7945,11685,13555,14424,7212,3606,1803,8612,4306,
                   2153,9749,12587,15028,7514,3757,9591,12442,6221,11783,13602,6801,12137,13717,14571,
                   15956,7978,3989,9707,12500,6250,3125,9275,12348,6174,3087,9254,4627,11048,5524,
                   2762,1381,8339,12904,6452,3226,1613,8455,12962,6481,11913,13669,14483,15976,7988,
                   3994,1997,8647,12994,6497,11921,13673,14485,15979,15636,7818,3909,9603,12512,6256,
                   3128,1564,782,391,8930,4465,10905,14189,14743,16106,8053,11675,13548,6774,3387,
                   9404,4702,2351,9910,4955,11148,5574,2787,10064,5032,2516,1258,629,8987,13228,
                   6614,3307,9300,4650,2325,9899,12660,6330,3165,9231,12326,6163,11816,5908,2954,
                   1477,8387,12864,6432,3216,1608,804,402,201,8773,13059,15264,7632,3816,1908,
                   954,477,8911,13126,6563,12016,6008,3004,1502,751,9046,4523,10996,5498,2749,
                   10111,12702,6351,11846,5923,10672,5336,2668,1334,667,9068,4534,2267,9804,4902,
                   2451,9960,4980,2490,1245,8271,12806,6403,11936,5968,2984,1492,746,373,8859,
                   13164,6582,3291,9292,4646,2323,9896,4948,2474,1237,8267,12804,6402,3201,9313,
                   12305,14889,16181,15803,15612,7806,3903,9662,4831,11086,5543,10482,5241,10269,13871,
                   14646,7323,11372,5686,2843,10156,5078,2539,9940,4970,2485,9979,12636,6318,3159,
                   9226,4613,11043,14256,7128,3564,1782,891,9116,4558,2279,9810,4905,11189,14331,
                   14812,7406,3703,9498,4749,11111,14226,7113,12229,13763,14528,7264,3632,1816,908,
                   454,227,8784,4392,2196,1098,549,9011,13240,6620,3310,1655,8474,4237,10855,
                   14098,7049,12261,13779,14536,7268,3634,1817,8621,13047,15194,7597,11511,13402,6701,
                   12087,13754,6877,12111,13702,6851,12096,6048,3024,1512,756,378,189,8831,13086,
                   6543,12006,6003,10648,5324,2662,1331,8376,4188,2094,1047,8234,4117,10795,14132,
                   7066,3533,9415,12354,6177,11825,13625,14525,15999,15646,7823,11622,5811,10616,5308,
                   2654,1327,8374,4187,10764,5382,2691,10080,5040,2520,1260,630,315,8892,4446,
                   2223,9846,4923,11196,5598,2799,10070,5035,11252,5626,2813,10079,12686,6343,11842,
                   5921,10673,14073,14685,16015,15718,7859,11640,5820,2910,1455,8438,4219,10780,5390,
                   2695,10082,5041,11257,14301,14799,16070,8035,11664,5832,2916,1458,729,9037,13191,
                   15330,7665,11481,13389,14343,15906,7953,11689,13557,14427,15884,7942,3971,9696,4848,
                   2424,1212,606,303,8886,4443,10892,5446,2723,10096,5048,2524,1262,631,8986,
                   4493,10983,14162,7081,12277,13787,14540,7270,3635,9528,4764,2382,1191,8306,4153,
                   10813,14143,14782,7391,11342,5671,10546,5273,10349,13847,14634,7317,11371,13332,6666,
                   3333,9379,12400,6200,3100,1550,775,9122,4561,10953,14149,14723,16096,8048,4024,
                   2012,1006,503,8922,4461,10903,14186,7093,12283,13788,6894,3447,9370,4685,11015,
                   14242,7121,12233,13765,14531,15936,7968,3984,1992,996,498,249,8797,13071,15270,
                   7635,11464,5732,2866,1433,8429,12887,15114,7557,11491,13392,6696,3348,1674,837,
                   9091,13280,6640,3320,1660,830,415,8942,4471,10906,5453,10375,13922,6961,12217,
                   13821,14559,15950,7975,11698,5849,10573,13959,14690,7345,11385,13341,14383,15926,7963,
                   11692,5846,2923,10132,5066,2533,9939,12616,6308,3154,1577,8501,12987,15228,7614,
                   3807,9550,4775,11122,5561,10493,13919,14606,7303,11362,5681,10553,14013,14719,16030,
                   8015,11654,5827,10560,5280,2640,1320,660,330,165,8819,13080,6540,3270,1635,
                   8464,4232,2116,1058,529,9001,13237,15355,16348,8174,4087,9690,4845,11095,14218,
                   7109,12227,13760,6880,3440,1720,860,430,215,8778,4389,10931,14200,7100,3550,
                   1775,8534,4267,10868,5434,2717,10095,12694,6347,11844,5922,2961,10217,12757,15051,
                   16196,8098,4049,9673,12485,14915,16128,8064,4032,2016,1008,504,252,126,63,
                   8766,4383,10926,5463,10378,5189,10243,13856,6928,3464,1732,866,433,8953,13149,
                   15247,16358,8179,11736,5868,2934,1467,8444,4222,2111,9790,4895,11182,5591,10442,
                   5221,10259,13864,6932,3466,1733,8515,12928,6464,3232,1616,808,404,202,101,
                   8723,13096,6548,3274,1637,8467,12968,6484,3242,1621,8459,12964,6482,3241,9333,
                   12315,14892,7446,3723,9572,4786,2393,9869,12647,14994,7497,11397,13411,14352,7176,
                   3588,1794,897,9185,13265,15305,16325,15811,15552,7776,3888,1944,972,486,243,
                   8792,4396,2198,1099,8196,4098,2049,9761,12593,15033,16253,15775,15598,7799,11546,
                   5773,10599,13970,6985,12165,13795,14544,7272,3636,1818,909,9191,13266,6633,11989,
                   13643,14468,7234,3617,9521,12473,14973,16159,15790,7895,11594,5797,10611,13976,6988,
                   3494,1747,8520,4260,2130,1065,8245,12859,15164,7582,3791,9542,4771,11120,5560,
                   2780,1390,695,9082,4541,11007,14174,7087,12278,6139,10716,5358,2679,10010,5005,
                   11239,14290,7145,12245,13771,14532,7266,3633,9529,12477,14975,16158,8079,11750,5875,
                   10584,5292,2646,1323,8372,4186,2093,9783,12602,6301,11887,13590,6795,12132,6066,
                   3033,10189,12743,15042,7521,11409,13417,14357,15915,15668,7834,3917,9607,12514,6257,
                   11801,13613,14519,15994,7997,11711,13566,6783,12062,6031,10726,5363,10328,5164,2582,
                   1291,8356,4178,2089,9781,12603,15036,7518,3759,9590,4795,11132,5566,2783,10062,
                   5031,11250,5625,10461,13903,14598,7299,11360,5680,2840,1420,710,355,8848,4424,
                   2212,1106,553,9013,13243,15356,7678,3839,9566,4783,11126,5563,10492,5246,2623,
                   10046,5023,11246,5623,10458,5229,10263,13866,6933,12203,13812,6906,3453,9375,12398,
                   6199,11834,5917,10671,14070,7035,12188,6094,3047,10194,5097,11221,14283,14788,7394,
                   3697,9497,12461,14967,16154,8077,11751,13522,6761,12053,13739,14580,7290,3645,9535,
                   12478,6239,11790,5895,10658,5329,10313,13829,14627,16048,8024,4012,2006,1003,9172,
                   4586,2293,9819,12556,6278,3139,9216,4608,2304,1152,576,288,144,72,36,
                   18,9,8741,13107,15288,7644,3822,1911,8602,4301,10823,14082,7041,12257,13777,
                   14537,15941,15619,15520,7760,3880,1940,970,485,8915,13128,6564,3282,1641,8469,
                   12971,15220,7610,3805,9551,12422,6211,11776,5888,2944,1472,736,368,184,92,
                   46,23,8746,4373,10923,14196,7098,3549,9423,12358,6179,11824,5912,2956,1478,
                   739,9040,4520,2260,1130,565,9019,13244,6622,3311,9302,4651,11060,5530,2765,
                   10055,12674,6337,11841,13569,14497,15985,15641,15533,15479,15386,7693,11559,13490,6745,
                   12045,13735,14578,7289,11293,13359,14390,7195,11308,5654,2827,10148,5074,2537,9941,
                   12619,14980,7490,3745,9585,12441,14957,16151,15786,7893,11595,13444,6722,3361,9393,
                   12409,14877,16175,15798,7899,11596,5798,2899,10120,5060,2530,1265,8281,12813,15143,
                   16306,8153,11725,13511,14402,7201,11313,13369,14397,15935,15678,7839,11630,5815,10618,
                   5309,10367,13854,6927,12198,6099,10696,5348,2674,1337,8381,12927,15134,7567,11494,
                   5747,10520,5260,2630,1315,8368,4184,2092,1046,523,8996,4498,2249,9797,12547,
                   15008,7504,3752,1876,938,469,8907,13124,6562,3281,9289,12293,14883,16176,8088,
                   4044,2022,1011,9176,4588,2294,1147,8220,4110,2055,9762,4881,11177,14325,14811,
                   16076,8038,4019,9720,4860,2430,1215,8318,4159,10814,5407,10414,5207,10250,5125,
                   10275,13872,6936,3468,1734,867,9104,4552,2276,1138,569,9021,13247,15358,7679,
                   11486,5743,10518,5259,10340,5170,2585,10029,12727,15098,7549,11423,13422,6711,12090,
                   6045,10735,14038,7019,12180,6090,3045,10195,12744,6372,3186,1593,8509,12991,15230,
                   7615,11518,5759,10526,5263,10342,5171,10296,5148,2574,1287,8354,4177,10761,14117,
                   14771,16120,8060,4030,2015,8654,4327,10834,5417,10421,13947,14620,7310,3655,9474,
                   4737,11105,14225,14825,16085,15691,15492,7746,3873,9649,12537,14941,16143,15782,7891,
                   11592,5796,2898,1449,8437,12891,15116,7558,3779,9536,4768,2384,1192,596,298,
                   149,8811,13076,6538,3269,9283,12288,6144,3072,1536,768,384,192,96,48,
                   24,12,6,3,8736,4368,2184,1092,546,273,8873,13173,15259,16364,8182,
                   4091,9692,4846,2423,9882,4941,11143,14306,7153,12249,13773,14535,15938,7969,11697,
                   13561,14429,15887,15654,7827,11624,5812,2906,1453,8439,12890,6445,11959,13690,6845,
                   12159,13726,6863,12102,6051,10736,5368,2684,1342,671,9070,4535,11002,5501,10399,
                   13934,6967,12218,6109,10703,14022,7011,12176,6088,3044,1522,761,9053,13199,15334,
                   7667,11480,5740,2870,1435,8428,4214,2107,9788,4894,2447,9958,4979,11160,5580,
                   2790,1395,8344,4172,2086,1043,8232,4116,2058,1029,8227,12848,6424,3212,1606,
                   803,9136,4568,2284,1142,571,9020,4510,2255,9798,4899,11184,5592,2796,1398,
                   699,9084,4542,2271,9806,4903,11186,5593,10445,13895,14594,7297,11361,13329,14377,
                   15925,15675,15548,7774,3887,9654,4827,11084,5542,2771,10056,5028,2514,1257,8277,
                   12811,15140,7570,3785,9541,12419,14944,7472,3736,1868,934,467,8904,4452,2226,
                   1113,8205,12839,15154,7577,11501,13399,14346,7173,11299,13360,6680,3340,1670,835,
                   9088,4544,2272,1136,568,284,142,71,8706,4353,10913,14193,14745,16109,15703,
                   15498,7749,11523,13472,6736,3368,1684,842,421,8947,13144,6572,3286,1643,8468,
                   4234,2117,9731,12576,6288,3144,1572,786,393,8933,13139,15240,7620,3810,1905,
                   8601,13037,15191,16266,8133,11715,13504,6752,3376,1688,844,422,211,8776,4388,
                   2194,1097,8197,12835,15152,7576,3788,1894,947,9208,4604,2302,1151,8222,4111,
                   10790,5395,10408,5204,2602,1301,8363,12916,6458,3229,9327,12310,6155,11812,5906,
                   2953,10213,12755,15048,7524,3762,1881,8589,13031,15186,7593,11509,13403,14348,7174,
                   3587,9504,4752,2376,1188,594,297,8885,13179,15260,7630,3815,9554,4777,11125,
                   14235,14828,7414,3707,9500,4750,2375,9858,4929,11137,14305,14801,16073,15685,15491,
                   15456,7728,3864,1932,966,483,8912,4456,2228,1114,557,9015,13242,6621,11983,
                   13638,6819,12144,6072,3036,1518,759,9050,4525,10999,14170,7085,12279,13786,6893,
                   12119,13706,6853,12099,13696,6848,3424,1712,856,428,214,107,8724,4362,2181,
                   9827,12560,6280,3140,1570,785,9129,13301,15323,16332,8166,4083,9688,4844,2422,
                   1211,8316,4158,2079,9774,4887,11178,5589,10443,13892,6946,3473,9449,12373,14859,
                   16164,8082,4041,9669,12483,14912,7456,3728,1864,932,466,233,8789,13067,15268,
                   7634,3817,9557,12427,14948,7474,3737,9581,12439,14954,7477,11451,13436,6718,3359,
                   9390,4695,11018,5509,10467,13904,6952,3476,1738,869,9107,13288,6644,3322,1661,
                   8479,12974,6487,11914,5957,10627,14048,7024,3512,1756,878,439,8954,4477,10911,
                   14190,7095,12282,6141,10719,14030,7015,12178,6089,10693,14019,14656,7328,3664,1832,
                   916,458,229,8787,13064,6532,3266,1633,8465,12969,15221,16283,15852,7926,3963,
                   9628,4814,2407,9874,4937,11141,14307,14800,7400,3700,1850,925,9199,13270,6635,
                   11988,5994,2997,10235,12764,6382,3191,9242,4621,11047,14258,7129,12237,13767,14530,
                   7265,11281,13353,14389,15931,15676,7838,3919,9606,4803,11072,5536,2768,1384,692,
                   346,173,8823,13082,6541,12007,13650,6825,12149,13723,14572,7286,3643,9532,4766,
                   2383,9862,4931,11136,5568,2784,1392,696,348,174,87,8714,4357,10915,14192,
                   7096,3548,1774,887,9114,4557,10951,14146,7073,12273,13785,14541,15943,15618,7809,
                   11617,13457,14441,15893,15659,15540,7770,3885,9655,12538,6269,11807,13614,6807,12138,
                   6069,10747,14044,7022,3511,9466,4733,11039,14254,7127,12234,6117,10707,14024,7012,
                   3506,1753,8525,12935,15202,7601,11513,13405,14351,15910,7955,11688,5844,2922,1461,
                   8443,12892,6446,3223,9322,4661,11067,14268,7134,3567,9430,4715,11028,5514,2757,
                   10051,12672,6336,3168,1584,792,396,198,99,8720,4360,2180,1090,545,9009,
                   13241,15357,16351,15822,7911,11602,5801,10613,13979,14700,7350,3675,9484,4742,2371,
                   9856,4928,2464,1232,616,308,154,77,8711,13090,6545,12009,13653,14475,15972,
                   7986,3993,9709,12503,14922,7461,11443,13432,6716,3358,1679,8550,4275,10872,5436,
                   2718,1359,8326,4163,10752,5376,2688,1344,672,336,168,84,42,21,8747,
                   13108,6554,3277,9287,12290,6145,11809,13617,14521,15997,15647,15534,7767,11530,5765,
                   10595,13968,6984,3492,1746,873,9109,13291,15316,7658,3829,9563,12428,6214,3107,
                   9264,4632,2316,1158,579,8960,4480,2240,1120,560,280,140,70,35,8752,
                   4376,2188,1094,547,9008,4504,2252,1126,563,9016,4508,2254,1127,8210,4105,
                   10789,14131,14776,7388,3694,1847,8634,4317,10831,14086,7043,12256,6128,3064,1532,
                   766,383,8862,4431,10886,5443,10368,5184,2592,1296,648,324,162,81,8713,
                   13093,15283,16376,8188,4094,2047,8670,4335,10838,5419,10420,5210,2605,10039,12730,
                   6365,11855,13574,6787,12128,6064,3032,1516,758,379,8860,4430,2215,9842,4921,
                   11197,14335,14814,7407,11350,5675,10548,5274,2637,9991,12706,6353,11849,13573,14499,
                   15984,7992,3996,1998,999,9170,4585,10965,14155,14724,7362,3681,9489,12457,14965,
                   16155,15788,7894,3947,9620,4810,2405,9875,12648,6324,3162,1581,8503,12986,6493,
                   11919,13670,6835,12152,6076,3038,1519,8406,4203,10772,5386,2693,10083,12688,6344,
                   3172,1586,793,9133,13303,15322,7661,11479,13386,6693,12083,13752,6876,3438,1719,
                   8570,4285,10879,14110,7055,12262,6131,10712,5356,2678,1339,8380,4190,2095,9782,
                   4891,11180,5590,2795,10068,5034,2517,9931,12612,6306,3153,9225,12325,14899,16184,
                   8092,4046,2023,8658,4329,10837,14091,14756,7378,3689,9493,12459,14964,7482,3741,
                   9583,12438,6219,11780,5890,2945,10209,12753,15049,16197,15747,15584,7792,3896,1948,
                   974,487,8914,4457,10901,14187,14740,7370,3685,9491,12456,6228,3114,1557,8491,
                   12980,6490,3245,9335,12314,6157,11815,13618,6809,12141,13719,14570,7285,11291,13356,
                   6678,3339,9380,4690,2345,9909,12667,15004,7502,3751,9586,4793,11133,14239,14830,
                   7415,11354,5677,10551,14010,7005,12175,13798,6899,12120,6060,3030,1515,8404,4202,
                   2101,9787,12604,6302,3151,9222,4611,11040,5520,2760,1380,690,345,8845,13159,
                   15250,7625,11461,13379,14336,7168,3584,1792,896,448,224,112,56,28,14,
                   7,8738,4369,10921,14197,14747,16108,8054,4027,9724,4862,2431,9886,4943,11142,
                   5571,10432,5216,2608,1304,652,326,163,8816,4408,2204,1102,551,9010,4505,
                   10989,14167,14730,7365,11331,13312,6656,3328,1664,832,416,208,104,52,26,
                   13,8743,13106,6553,12013,13655,14474,7237,11267,13344,6672,3336,1668,834,417,
                   8945,13145,15245,16359,15826,7913,11605,13451,14436,7218,3609,9517,12471,14970,7485,
                   11455,13438,6719,12094,6047,10734,5367,10330,5165,10295,13882,6941,12207,13814,6907,
                   12124,6062,3031,10186,5093,11219,14280,7140,3570,1785,8541,12943,15206,7603,11512,
                   5756,2878,1439,8430,4215,10778,5389,10407,13938,6969,12221,13823,14558,7279,11286,
                   5643,10532,5266,2633,9989,12707,15088,7544,3772,1886,943,9206,4603,10972,5486,
                   2743,10106,5053,11263,14302,7151,12246,6123,10708,5354,2677,10011,12716,6358,3179,
                   9236,4618,2309,9891,12656,6328,3164,1582,791,9130,4565,10955,14148,7074,3537,
                   9417,12357,14851,16160,8080,4040,2020,1010,505,8925,13135,15238,7619,11456,5728,
                   2864,1432,716,358,179,8824,4412,2206,1103,8198,4099,10784,5392,2696,1348,
                   674,337,8841,13157,15251,16360,8180,4090,2045,8671,13006,6503,11922,5961,10629,
                   14051,14672,7336,3668,1834,917,9195,13268,6634,3317,9307,12300,6150,3075,9248,
                   4624,2312,1156,578,289,8881,13177,15261,16367,15830,7915,11604,5802,2901,10123,
                   12772,6386,3193,9245,12335,14902,7451,11436,5718,2859,10164,5082,2541,9943,12618,
                   6309,11891,13592,6796,3398,1699,8560,4280,2140,1070,535,9002,4501,10987,14164,
                   7082,3541,9419,12356,6178,3089,9257,12341,14907,16188,8094,4047,9670,4835,11088,
                   5544,2772,1386,693,9083,13212,6606,3303,9298,4649,11061,14267,14844,7422,3711,
                   9502,4751,11110,5555,10488,5244,2622,1311,8366,4183,10762,5381,10403,13936,6968,
                   3484,1742,871,9106,4553,10949,14147,14720,7360,3680,1840,920,460,230,115,
                   8728,4364,2182,1091,8192,4096,2048,1024,512,256,128,64,32,16,8,
                   4,2,1);
constant powernum : numarray := (1,2,4,8,16,32,64,128,256,512,1024,2048,4096,8192,1091,2182,
                   4364,8728,115,230,460,920,1840,3680,7360,14720,14147,10949,4553,9106,871,
                   1742,3484,6968,13936,10403,5381,10762,4183,8366,1311,2622,5244,10488,5555,11110,
                   4751,9502,3711,7422,14844,14267,11061,4649,9298,3303,6606,13212,9083,693,1386,
                   2772,5544,11088,4835,9670,4047,8094,16188,14907,12341,9257,3089,6178,12356,9419,
                   3541,7082,14164,10987,4501,9002,535,1070,2140,4280,8560,1699,3398,6796,13592,
                   11891,6309,12618,9943,2541,5082,10164,2859,5718,11436,7451,14902,12335,9245,3193,
                   6386,12772,10123,2901,5802,11604,7915,15830,16367,15261,13177,8881,289,578,1156,
                   2312,4624,9248,3075,6150,12300,9307,3317,6634,13268,9195,917,1834,3668,7336,
                   14672,14051,10629,5961,11922,6503,13006,8671,2045,4090,8180,16360,15251,13157,8841,
                   337,674,1348,2696,5392,10784,4099,8198,1103,2206,4412,8824,179,358,716,
                   1432,2864,5728,11456,7619,15238,13135,8925,505,1010,2020,4040,8080,16160,14851,
                   12357,9417,3537,7074,14148,10955,4565,9130,791,1582,3164,6328,12656,9891,2309,
                   4618,9236,3179,6358,12716,10011,2677,5354,10708,6123,12246,7151,14302,11263,5053,
                   10106,2743,5486,10972,4603,9206,943,1886,3772,7544,15088,12707,9989,2633,5266,
                   10532,5643,11286,7279,14558,13823,12221,6969,13938,10407,5389,10778,4215,8430,1439,
                   2878,5756,11512,7603,15206,12943,8541,1785,3570,7140,14280,11219,5093,10186,3031,
                   6062,12124,6907,13814,12207,6941,13882,10295,5165,10330,5367,10734,6047,12094,6719,
                   13438,11455,7485,14970,12471,9517,3609,7218,14436,13451,11605,7913,15826,16359,15245,
                   13145,8945,417,834,1668,3336,6672,13344,11267,7237,14474,13655,12013,6553,13106,
                   8743,13,26,52,104,208,416,832,1664,3328,6656,13312,11331,7365,14730,
                   14167,10989,4505,9010,551,1102,2204,4408,8816,163,326,652,1304,2608,5216,
                   10432,5571,11142,4943,9886,2431,4862,9724,4027,8054,16108,14747,14197,10921,4369,
                   8738,7,14,28,56,112,224,448,896,1792,3584,7168,14336,13379,11461,
                   7625,15250,13159,8845,345,690,1380,2760,5520,11040,4611,9222,3151,6302,12604,
                   9787,2101,4202,8404,1515,3030,6060,12120,6899,13798,12175,7005,14010,10551,5677,
                   11354,7415,14830,14239,11133,4793,9586,3751,7502,15004,12667,9909,2345,4690,9380,
                   3339,6678,13356,11291,7285,14570,13719,12141,6809,13618,11815,6157,12314,9335,3245,
                   6490,12980,8491,1557,3114,6228,12456,9491,3685,7370,14740,14187,10901,4457,8914,
                   487,974,1948,3896,7792,15584,15747,16197,15049,12753,10209,2945,5890,11780,6219,
                   12438,9583,3741,7482,14964,12459,9493,3689,7378,14756,14091,10837,4329,8658,2023,
                   4046,8092,16184,14899,12325,9225,3153,6306,12612,9931,2517,5034,10068,2795,5590,
                   11180,4891,9782,2095,4190,8380,1339,2678,5356,10712,6131,12262,7055,14110,10879,
                   4285,8570,1719,3438,6876,13752,12083,6693,13386,11479,7661,15322,13303,9133,793,
                   1586,3172,6344,12688,10083,2693,5386,10772,4203,8406,1519,3038,6076,12152,6835,
                   13670,11919,6493,12986,8503,1581,3162,6324,12648,9875,2405,4810,9620,3947,7894,
                   15788,16155,14965,12457,9489,3681,7362,14724,14155,10965,4585,9170,999,1998,3996,
                   7992,15984,14499,13573,11849,6353,12706,9991,2637,5274,10548,5675,11350,7407,14814,
                   14335,11197,4921,9842,2215,4430,8860,379,758,1516,3032,6064,12128,6787,13574,
                   11855,6365,12730,10039,2605,5210,10420,5419,10838,4335,8670,2047,4094,8188,16376,
                   15283,13093,8713,81,162,324,648,1296,2592,5184,10368,5443,10886,4431,8862,
                   383,766,1532,3064,6128,12256,7043,14086,10831,4317,8634,1847,3694,7388,14776,
                   14131,10789,4105,8210,1127,2254,4508,9016,563,1126,2252,4504,9008,547,1094,
                   2188,4376,8752,35,70,140,280,560,1120,2240,4480,8960,579,1158,2316,
                   4632,9264,3107,6214,12428,9563,3829,7658,15316,13291,9109,873,1746,3492,6984,
                   13968,10595,5765,11530,7767,15534,15647,15997,14521,13617,11809,6145,12290,9287,3277,
                   6554,13108,8747,21,42,84,168,336,672,1344,2688,5376,10752,4163,8326,
                   1359,2718,5436,10872,4275,8550,1679,3358,6716,13432,11443,7461,14922,12503,9709,
                   3993,7986,15972,14475,13653,12009,6545,13090,8711,77,154,308,616,1232,2464,
                   4928,9856,2371,4742,9484,3675,7350,14700,13979,10613,5801,11602,7911,15822,16351,
                   15357,13241,9009,545,1090,2180,4360,8720,99,198,396,792,1584,3168,6336,
                   12672,10051,2757,5514,11028,4715,9430,3567,7134,14268,11067,4661,9322,3223,6446,
                   12892,8443,1461,2922,5844,11688,7955,15910,14351,13405,11513,7601,15202,12935,8525,
                   1753,3506,7012,14024,10707,6117,12234,7127,14254,11039,4733,9466,3511,7022,14044,
                   10747,6069,12138,6807,13614,11807,6269,12538,9655,3885,7770,15540,15659,15893,14441,
                   13457,11617,7809,15618,15943,14541,13785,12273,7073,14146,10951,4557,9114,887,1774,
                   3548,7096,14192,10915,4357,8714,87,174,348,696,1392,2784,5568,11136,4931,
                   9862,2383,4766,9532,3643,7286,14572,13723,12149,6825,13650,12007,6541,13082,8823,
                   173,346,692,1384,2768,5536,11072,4803,9606,3919,7838,15676,15931,14389,13353,
                   11281,7265,14530,13767,12237,7129,14258,11047,4621,9242,3191,6382,12764,10235,2997,
                   5994,11988,6635,13270,9199,925,1850,3700,7400,14800,14307,11141,4937,9874,2407,
                   4814,9628,3963,7926,15852,16283,15221,12969,8465,1633,3266,6532,13064,8787,229,
                   458,916,1832,3664,7328,14656,14019,10693,6089,12178,7015,14030,10719,6141,12282,
                   7095,14190,10911,4477,8954,439,878,1756,3512,7024,14048,10627,5957,11914,6487,
                   12974,8479,1661,3322,6644,13288,9107,869,1738,3476,6952,13904,10467,5509,11018,
                   4695,9390,3359,6718,13436,11451,7477,14954,12439,9581,3737,7474,14948,12427,9557,
                   3817,7634,15268,13067,8789,233,466,932,1864,3728,7456,14912,12483,9669,4041,
                   8082,16164,14859,12373,9449,3473,6946,13892,10443,5589,11178,4887,9774,2079,4158,
                   8316,1211,2422,4844,9688,4083,8166,16332,15323,13301,9129,785,1570,3140,6280,
                   12560,9827,2181,4362,8724,107,214,428,856,1712,3424,6848,13696,12099,6853,
                   13706,12119,6893,13786,12279,7085,14170,10999,4525,9050,759,1518,3036,6072,12144,
                   6819,13638,11983,6621,13242,9015,557,1114,2228,4456,8912,483,966,1932,3864,
                   7728,15456,15491,15685,16073,14801,14305,11137,4929,9858,2375,4750,9500,3707,7414,
                   14828,14235,11125,4777,9554,3815,7630,15260,13179,8885,297,594,1188,2376,4752,
                   9504,3587,7174,14348,13403,11509,7593,15186,13031,8589,1881,3762,7524,15048,12755,
                   10213,2953,5906,11812,6155,12310,9327,3229,6458,12916,8363,1301,2602,5204,10408,
                   5395,10790,4111,8222,1151,2302,4604,9208,947,1894,3788,7576,15152,12835,8197,
                   1097,2194,4388,8776,211,422,844,1688,3376,6752,13504,11715,8133,16266,15191,
                   13037,8601,1905,3810,7620,15240,13139,8933,393,786,1572,3144,6288,12576,9731,
                   2117,4234,8468,1643,3286,6572,13144,8947,421,842,1684,3368,6736,13472,11523,
                   7749,15498,15703,16109,14745,14193,10913,4353,8706,71,142,284,568,1136,2272,
                   4544,9088,835,1670,3340,6680,13360,11299,7173,14346,13399,11501,7577,15154,12839,
                   8205,1113,2226,4452,8904,467,934,1868,3736,7472,14944,12419,9541,3785,7570,
                   15140,12811,8277,1257,2514,5028,10056,2771,5542,11084,4827,9654,3887,7774,15548,
                   15675,15925,14377,13329,11361,7297,14594,13895,10445,5593,11186,4903,9806,2271,4542,
                   9084,699,1398,2796,5592,11184,4899,9798,2255,4510,9020,571,1142,2284,4568,
                   9136,803,1606,3212,6424,12848,8227,1029,2058,4116,8232,1043,2086,4172,8344,
                   1395,2790,5580,11160,4979,9958,2447,4894,9788,2107,4214,8428,1435,2870,5740,
                   11480,7667,15334,13199,9053,761,1522,3044,6088,12176,7011,14022,10703,6109,12218,
                   6967,13934,10399,5501,11002,4535,9070,671,1342,2684,5368,10736,6051,12102,6863,
                   13726,12159,6845,13690,11959,6445,12890,8439,1453,2906,5812,11624,7827,15654,15887,
                   14429,13561,11697,7969,15938,14535,13773,12249,7153,14306,11143,4941,9882,2423,4846,
                   9692,4091,8182,16364,15259,13173,8873,273,546,1092,2184,4368,8736,3,6,
                   12,24,48,96,192,384,768,1536,3072,6144,12288,9283,3269,6538,13076,
                   8811,149,298,596,1192,2384,4768,9536,3779,7558,15116,12891,8437,1449,2898,
                   5796,11592,7891,15782,16143,14941,12537,9649,3873,7746,15492,15691,16085,14825,14225,
                   11105,4737,9474,3655,7310,14620,13947,10421,5417,10834,4327,8654,2015,4030,8060,
                   16120,14771,14117,10761,4177,8354,1287,2574,5148,10296,5171,10342,5263,10526,5759,
                   11518,7615,15230,12991,8509,1593,3186,6372,12744,10195,3045,6090,12180,7019,14038,
                   10735,6045,12090,6711,13422,11423,7549,15098,12727,10029,2585,5170,10340,5259,10518,
                   5743,11486,7679,15358,13247,9021,569,1138,2276,4552,9104,867,1734,3468,6936,
                   13872,10275,5125,10250,5207,10414,5407,10814,4159,8318,1215,2430,4860,9720,4019,
                   8038,16076,14811,14325,11177,4881,9762,2055,4110,8220,1147,2294,4588,9176,1011,
                   2022,4044,8088,16176,14883,12293,9289,3281,6562,13124,8907,469,938,1876,3752,
                   7504,15008,12547,9797,2249,4498,8996,523,1046,2092,4184,8368,1315,2630,5260,
                   10520,5747,11494,7567,15134,12927,8381,1337,2674,5348,10696,6099,12198,6927,13854,
                   10367,5309,10618,5815,11630,7839,15678,15935,14397,13369,11313,7201,14402,13511,11725,
                   8153,16306,15143,12813,8281,1265,2530,5060,10120,2899,5798,11596,7899,15798,16175,
                   14877,12409,9393,3361,6722,13444,11595,7893,15786,16151,14957,12441,9585,3745,7490,
                   14980,12619,9941,2537,5074,10148,2827,5654,11308,7195,14390,13359,11293,7289,14578,
                   13735,12045,6745,13490,11559,7693,15386,15479,15533,15641,15985,14497,13569,11841,6337,
                   12674,10055,2765,5530,11060,4651,9302,3311,6622,13244,9019,565,1130,2260,4520,
                   9040,739,1478,2956,5912,11824,6179,12358,9423,3549,7098,14196,10923,4373,8746,
                   23,46,92,184,368,736,1472,2944,5888,11776,6211,12422,9551,3805,7610,
                   15220,12971,8469,1641,3282,6564,13128,8915,485,970,1940,3880,7760,15520,15619,
                   15941,14537,13777,12257,7041,14082,10823,4301,8602,1911,3822,7644,15288,13107,8741,
                   9,18,36,72,144,288,576,1152,2304,4608,9216,3139,6278,12556,9819,
                   2293,4586,9172,1003,2006,4012,8024,16048,14627,13829,10313,5329,10658,5895,11790,
                   6239,12478,9535,3645,7290,14580,13739,12053,6761,13522,11751,8077,16154,14967,12461,
                   9497,3697,7394,14788,14283,11221,5097,10194,3047,6094,12188,7035,14070,10671,5917,
                   11834,6199,12398,9375,3453,6906,13812,12203,6933,13866,10263,5229,10458,5623,11246,
                   5023,10046,2623,5246,10492,5563,11126,4783,9566,3839,7678,15356,13243,9013,553,
                   1106,2212,4424,8848,355,710,1420,2840,5680,11360,7299,14598,13903,10461,5625,
                   11250,5031,10062,2783,5566,11132,4795,9590,3759,7518,15036,12603,9781,2089,4178,
                   8356,1291,2582,5164,10328,5363,10726,6031,12062,6783,13566,11711,7997,15994,14519,
                   13613,11801,6257,12514,9607,3917,7834,15668,15915,14357,13417,11409,7521,15042,12743,
                   10189,3033,6066,12132,6795,13590,11887,6301,12602,9783,2093,4186,8372,1323,2646,
                   5292,10584,5875,11750,8079,16158,14975,12477,9529,3633,7266,14532,13771,12245,7145,
                   14290,11239,5005,10010,2679,5358,10716,6139,12278,7087,14174,11007,4541,9082,695,
                   1390,2780,5560,11120,4771,9542,3791,7582,15164,12859,8245,1065,2130,4260,8520,
                   1747,3494,6988,13976,10611,5797,11594,7895,15790,16159,14973,12473,9521,3617,7234,
                   14468,13643,11989,6633,13266,9191,909,1818,3636,7272,14544,13795,12165,6985,13970,
                   10599,5773,11546,7799,15598,15775,16253,15033,12593,9761,2049,4098,8196,1099,2198,
                   4396,8792,243,486,972,1944,3888,7776,15552,15811,16325,15305,13265,9185,897,
                   1794,3588,7176,14352,13411,11397,7497,14994,12647,9869,2393,4786,9572,3723,7446,
                   14892,12315,9333,3241,6482,12964,8459,1621,3242,6484,12968,8467,1637,3274,6548,
                   13096,8723,101,202,404,808,1616,3232,6464,12928,8515,1733,3466,6932,13864,
                   10259,5221,10442,5591,11182,4895,9790,2111,4222,8444,1467,2934,5868,11736,8179,
                   16358,15247,13149,8953,433,866,1732,3464,6928,13856,10243,5189,10378,5463,10926,
                   4383,8766,63,126,252,504,1008,2016,4032,8064,16128,14915,12485,9673,4049,
                   8098,16196,15051,12757,10217,2961,5922,11844,6347,12694,10095,2717,5434,10868,4267,
                   8534,1775,3550,7100,14200,10931,4389,8778,215,430,860,1720,3440,6880,13760,
                   12227,7109,14218,11095,4845,9690,4087,8174,16348,15355,13237,9001,529,1058,2116,
                   4232,8464,1635,3270,6540,13080,8819,165,330,660,1320,2640,5280,10560,5827,
                   11654,8015,16030,14719,14013,10553,5681,11362,7303,14606,13919,10493,5561,11122,4775,
                   9550,3807,7614,15228,12987,8501,1577,3154,6308,12616,9939,2533,5066,10132,2923,
                   5846,11692,7963,15926,14383,13341,11385,7345,14690,13959,10573,5849,11698,7975,15950,
                   14559,13821,12217,6961,13922,10375,5453,10906,4471,8942,415,830,1660,3320,6640,
                   13280,9091,837,1674,3348,6696,13392,11491,7557,15114,12887,8429,1433,2866,5732,
                   11464,7635,15270,13071,8797,249,498,996,1992,3984,7968,15936,14531,13765,12233,
                   7121,14242,11015,4685,9370,3447,6894,13788,12283,7093,14186,10903,4461,8922,503,
                   1006,2012,4024,8048,16096,14723,14149,10953,4561,9122,775,1550,3100,6200,12400,
                   9379,3333,6666,13332,11371,7317,14634,13847,10349,5273,10546,5671,11342,7391,14782,
                   14143,10813,4153,8306,1191,2382,4764,9528,3635,7270,14540,13787,12277,7081,14162,
                   10983,4493,8986,631,1262,2524,5048,10096,2723,5446,10892,4443,8886,303,606,
                   1212,2424,4848,9696,3971,7942,15884,14427,13557,11689,7953,15906,14343,13389,11481,
                   7665,15330,13191,9037,729,1458,2916,5832,11664,8035,16070,14799,14301,11257,5041,
                   10082,2695,5390,10780,4219,8438,1455,2910,5820,11640,7859,15718,16015,14685,14073,
                   10673,5921,11842,6343,12686,10079,2813,5626,11252,5035,10070,2799,5598,11196,4923,
                   9846,2223,4446,8892,315,630,1260,2520,5040,10080,2691,5382,10764,4187,8374,
                   1327,2654,5308,10616,5811,11622,7823,15646,15999,14525,13625,11825,6177,12354,9415,
                   3533,7066,14132,10795,4117,8234,1047,2094,4188,8376,1331,2662,5324,10648,6003,
                   12006,6543,13086,8831,189,378,756,1512,3024,6048,12096,6851,13702,12111,6877,
                   13754,12087,6701,13402,11511,7597,15194,13047,8621,1817,3634,7268,14536,13779,12261,
                   7049,14098,10855,4237,8474,1655,3310,6620,13240,9011,549,1098,2196,4392,8784,
                   227,454,908,1816,3632,7264,14528,13763,12229,7113,14226,11111,4749,9498,3703,
                   7406,14812,14331,11189,4905,9810,2279,4558,9116,891,1782,3564,7128,14256,11043,
                   4613,9226,3159,6318,12636,9979,2485,4970,9940,2539,5078,10156,2843,5686,11372,
                   7323,14646,13871,10269,5241,10482,5543,11086,4831,9662,3903,7806,15612,15803,16181,
                   14889,12305,9313,3201,6402,12804,8267,1237,2474,4948,9896,2323,4646,9292,3291,
                   6582,13164,8859,373,746,1492,2984,5968,11936,6403,12806,8271,1245,2490,4980,
                   9960,2451,4902,9804,2267,4534,9068,667,1334,2668,5336,10672,5923,11846,6351,
                   12702,10111,2749,5498,10996,4523,9046,751,1502,3004,6008,12016,6563,13126,8911,
                   477,954,1908,3816,7632,15264,13059,8773,201,402,804,1608,3216,6432,12864,
                   8387,1477,2954,5908,11816,6163,12326,9231,3165,6330,12660,9899,2325,4650,9300,
                   3307,6614,13228,8987,629,1258,2516,5032,10064,2787,5574,11148,4955,9910,2351,
                   4702,9404,3387,6774,13548,11675,8053,16106,14743,14189,10905,4465,8930,391,782,
                   1564,3128,6256,12512,9603,3909,7818,15636,15979,14485,13673,11921,6497,12994,8647,
                   1997,3994,7988,15976,14483,13669,11913,6481,12962,8455,1613,3226,6452,12904,8339,
                   1381,2762,5524,11048,4627,9254,3087,6174,12348,9275,3125,6250,12500,9707,3989,
                   7978,15956,14571,13717,12137,6801,13602,11783,6221,12442,9591,3757,7514,15028,12587,
                   9749,2153,4306,8612,1803,3606,7212,14424,13555,11685,7945,15890,14439,13453,11609,
                   7921,15842,16263,15181,13017,8689,1953,3906,7812,15624,15955,14565,13705,12113,6881,
                   13762,12231,7117,14234,11127,4781,9562,3831,7662,15324,13307,9141,809,1618,3236,
                   6472,12944,8547,1669,3338,6676,13352,11283,7269,14538,13783,12269,7065,14130,10791,
                   4109,8218,1143,2286,4572,9144,819,1638,3276,6552,13104,8739,5,10,20,
                   40,80,160,320,640,1280,2560,5120,10240,5187,10374,5455,10910,4479,8958,
                   447,894,1788,3576,7152,14304,11139,4933,9866,2391,4782,9564,3835,7670,15340,
                   13211,9077,681,1362,2724,5448,10896,4451,8902,463,926,1852,3704,7408,14816,
                   14211,11077,4809,9618,3943,7886,15772,16251,15029,12585,9745,2145,4290,8580,1867,
                   3734,7468,14936,12531,9637,3849,7698,15396,15371,15445,15593,15761,16225,14977,12609,
                   9921,2497,4994,9988,2635,5270,10540,5659,11318,7215,14430,13567,11709,7993,15986,
                   14503,13581,11865,6385,12770,10119,2893,5786,11572,7723,15446,15599,15773,16249,15025,
                   12577,9729,2113,4226,8452,1611,3222,6444,12888,8435,1445,2890,5780,11560,7699,
                   15398,15375,15453,15609,15793,16161,14849,12353,9409,3521,7042,14084,10827,4309,8618,
                   1815,3630,7260,14520,13619,11813,6153,12306,9319,3213,6426,12852,8235,1045,2090,
                   4180,8360,1299,2598,5196,10392,5491,10982,4495,8990,639,1278,2556,5112,10224,
                   2979,5958,11916,6491,12982,8495,1565,3130,6260,12520,9619,3941,7882,15764,16235,
                   14997,12649,9873,2401,4802,9604,3915,7830,15660,15899,14453,13481,11537,7777,15554,
                   15815,16333,15321,13297,9121,769,1538,3076,6152,12304,9315,3205,6410,12820,8299,
                   1173,2346,4692,9384,3347,6694,13388,11483,7669,15338,13207,9069,665,1330,2660,
                   5320,10640,5987,11974,6607,13214,9087,701,1402,2804,5608,11216,5091,10182,3023,
                   6046,12092,6715,13430,11439,7453,14906,12343,9261,3097,6194,12388,9355,3413,6826,
                   13652,12011,6549,13098,8727,109,218,436,872,1744,3488,6976,13952,10563,5829,
                   11658,8023,16046,14623,13949,10425,5425,10850,4231,8462,1631,3262,6524,13048,8627,
                   1829,3658,7316,14632,13843,10341,5257,10514,5735,11470,7647,15294,13119,8765,57,
                   114,228,456,912,1824,3648,7296,14592,13891,10437,5577,11154,4967,9934,2527,
                   5054,10108,2747,5494,10988,4507,9014,559,1118,2236,4472,8944,419,838,1676,
                   3352,6704,13408,11395,7493,14986,12631,9965,2457,4914,9828,2187,4374,8748,27,
                   54,108,216,432,864,1728,3456,6912,13824,10307,5317,10634,5975,11950,6431,
                   12862,8255,1085,2170,4340,8680,1939,3878,7756,15512,15731,16037,14601,13905,10465,
                   5505,11010,4679,9358,3423,6846,13692,11963,6453,12906,8343,1389,2778,5556,11112,
                   4755,9510,3599,7198,14396,13371,11317,7209,14418,13543,11661,8025,16050,14631,13837,
                   10329,5361,10722,6023,12046,6751,13502,11583,7741,15482,15543,15661,15897,14449,13473,
                   11521,7745,15490,15687,16077,14809,14321,11169,4865,9730,2119,4238,8476,1659,3318,
                   6636,13272,9203,933,1866,3732,7464,14928,12515,9605,3913,7826,15652,15883,14421,
                   13545,11665,8033,16066,14791,14285,11225,5105,10210,2951,5902,11804,6267,12534,9647,
                   3869,7738,15476,15531,15637,15977,14481,13665,11905,6465,12930,8519,1741,3482,6964,
                   13928,10387,5477,10954,4567,9134,799,1598,3196,6392,12784,10147,2821,5642,11284,
                   7275,14550,13807,12189,7033,14066,10663,5901,11802,6263,12526,9631,3965,7930,15860,
                   16299,15125,12905,8337,1377,2754,5508,11016,4691,9382,3343,6686,13372,11323,7221,
                   14442,13463,11629,7833,15666,15911,14349,13401,11505,7585,15170,12999,8653,2009,4018,
                   8036,16072,14803,14309,11145,4945,9890,2311,4622,9244,3195,6390,12780,10139,2933,
                   5866,11732,8171,16342,15343,13213,9081,689,1378,2756,5512,11024,4707,9414,3535,
                   7070,14140,10811,4149,8298,1175,2350,4700,9400,3379,6758,13516,11739,8181,16362,
                   15255,13165,8857,369,738,1476,2952,5904,11808,6147,12294,9295,3293,6586,13172,
                   8875,277,554,1108,2216,4432,8864,259,518,1036,2072,4144,8288,1155,2310,
                   4620,9240,3187,6374,12748,10203,3061,6122,12244,7147,14294,11247,5021,10042,2615,
                   5230,10460,5627,11254,5039,10078,2815,5630,11260,5051,10102,2735,5470,10940,4411,
                   8822,175,350,700,1400,2800,5600,11200,5059,10118,2895,5790,11580,7739,15478,
                   15535,15645,15993,14513,13601,11777,6209,12418,9543,3789,7578,15156,12843,8213,1129,
                   2258,4516,9032,723,1446,2892,5784,11568,7715,15430,15567,15837,16377,15281,13089,
                   8705,65,130,260,520,1040,2080,4160,8320,1347,2694,5388,10776,4211,8422,
                   1423,2846,5692,11384,7347,14694,13967,10589,5881,11762,8103,16206,15071,12797,10169,
                   2865,5730,11460,7627,15254,13167,8861,377,754,1508,3016,6032,12064,6659,13318,
                   11343,7389,14778,14135,10797,4121,8242,1063,2126,4252,8504,1587,3174,6348,12696,
                   10099,2725,5450,10900,4459,8918,495,990,1980,3960,7920,15840,16259,15173,13001,
                   8657,2017,4034,8068,16136,14931,12517,9609,3921,7842,15684,16075,14805,14313,11153,
                   4961,9922,2503,5006,10012,2683,5366,10732,6043,12086,6703,13406,11519,7613,15226,
                   12983,8493,1561,3122,6244,12488,9683,4069,8138,16276,15211,12949,8553,1681,3362,
                   6724,13448,11603,7909,15818,16343,15341,13209,9073,673,1346,2692,5384,10768,4195,
                   8390,1487,2974,5948,11896,6323,12646,9871,2397,4794,9588,3755,7510,15020,12571,
                   9845,2217,4434,8868,267,534,1068,2136,4272,8544,1667,3334,6668,13336,11379,
                   7333,14666,14039,10733,6041,12082,6695,13390,11487,7677,15354,13239,9005,537,1074,
                   2148,4296,8592,1891,3782,7564,15128,12915,8357,1289,2578,5156,10312,5331,10662,
                   5903,11806,6271,12542,9663,3901,7802,15604,15787,16149,14953,12433,9569,3713,7426,
                   14852,12363,9429,3561,7122,14244,11019,4693,9386,3351,6702,13404,11515,7605,15210,
                   12951,8557,1689,3378,6756,13512,11731,8165,16330,15319,13293,9113,881,1762,3524,
                   7048,14096,10851,4229,8458,1623,3246,6492,12984,8499,1573,3146,6292,12584,9747,
                   2149,4298,8596,1899,3798,7596,15192,13043,8613,1801,3602,7204,14408,13523,11749,
                   8073,16146,14951,12429,9561,3825,7650,15300,13259,9173,1001,2002,4004,8008,16016,
                   14691,13957,10569,5841,11682,7943,15886,14431,13565,11705,7985,15970,14471,13645,11993,
                   6641,13282,9095,845,1690,3380,6760,13520,11747,8069,16138,14935,12525,9625,3953,
                   7906,15812,16331,15317,13289,9105,865,1730,3460,6920,13840,10339,5253,10506,5719,
                   11438,7455,14910,12351,9277,3129,6258,12516,9611,3925,7850,15700,16107,14741,14185,
                   10897,4449,8898,455,910,1820,3640,7280,14560,13699,12101,6857,13714,12135,6797,
                   13594,11895,6317,12634,9975,2477,4954,9908,2347,4694,9388,3355,6710,13420,11419,
                   7541,15082,12695,10093,2713,5426,10852,4235,8470,1647,3294,6588,13176,8883,293,
                   586,1172,2344,4688,9376,3331,6662,13324,11355,7413,14826,14231,11117,4761,9522,
                   3623,7246,14492,13691,11957,6441,12882,8423,1421,2842,5684,11368,7315,14630,13839,
                   10333,5369,10738,6055,12110,6879,13758,12095,6717,13434,11447,7469,14938,12535,9645,
                   3865,7730,15460,15499,15701,16105,14737,14177,10881,4417,8834,327,654,1308,2616,
                   5232,10464,5507,11014,4687,9374,3455,6910,13820,12219,6965,13930,10391,5485,10970,
                   4599,9198,927,1854,3708,7416,14832,14243,11013,4681,9362,3431,6862,13724,12155,
                   6837,13674,11927,6509,13018,8695,1965,3930,7860,15720,16019,14693,13961,10577,5857,
                   11714,8135,16270,15199,13053,8633,1841,3682,7364,14728,14163,10981,4489,8978,615,
                   1230,2460,4920,9840,2211,4422,8844,347,694,1388,2776,5552,11104,4739,9478,
                   3663,7326,14652,13883,10293,5161,10322,5351,10702,6111,12222,6975,13950,10431,5437,
                   10874,4279,8558,1695,3390,6780,13560,11699,7973,15946,14551,13805,12185,7025,14050,
                   10631,5965,11930,6519,13038,8607,1917,3834,7668,15336,13203,9061,649,1298,2596,
                   5192,10384,5475,10950,4559,9118,895,1790,3580,7160,14320,11171,4869,9738,2135,
                   4270,8540,1787,3574,7148,14296,11251,5029,10058,2775,5550,11100,4859,9718,4015,
                   8030,16060,14651,13877,10281,5137,10274,5127,10254,5215,10430,5439,10878,4287,8574,
                   1727,3454,6908,13816,12211,6949,13898,10455,5613,11226,5111,10222,2975,5950,11900,
                   6331,12662,9903,2333,4666,9332,3243,6486,12972,8475,1653,3306,6612,13224,8979,
                   613,1226,2452,4904,9808,2275,4550,9100,859,1718,3436,6872,13744,12067,6661,
                   13322,11351,7405,14810,14327,11181,4889,9778,2087,4174,8348,1403,2806,5612,11224,
                   5107,10214,2959,5918,11836,6203,12406,9391,3357,6714,13428,11435,7445,14890,12311,
                   9325,3225,6450,12900,8331,1365,2730,5460,10920,4371,8742,15,30,60,120,
                   240,480,960,1920,3840,7680,15360,15427,15557,15817,16337,15329,13185,9025,705,
                   1410,2820,5640,11280,7267,14534,13775,12253,7161,14322,11175,4877,9754,2167,4334,
                   8668,2043,4086,8172,16344,15347,13221,8969,593,1186,2372,4744,9488,3683,7366,
                   14732,14171,10997,4521,9042,743,1486,2972,5944,11888,6307,12614,9935,2525,5050,
                   10100,2731,5462,10924,4379,8758,47,94,188,376,752,1504,3008,6016,12032,
                   6723,13446,11599,7901,15802,16183,14893,12313,9329,3233,6466,12932,8523,1749,3498,
                   6996,13992,10515,5733,11466,7639,15278,13087,8829,185,370,740,1480,2960,5920,
                   11840,6339,12678,10063,2781,5562,11124,4779,9558,3823,7646,15292,13115,8757,41,
                   82,164,328,656,1312,2624,5248,10496,5699,11398,7503,15006,12671,9917,2361,
                   4722,9444,3467,6934,13868,10267,5237,10474,5527,11054,4639,9278,3135,6270,12540,
                   9659,3893,7786,15572,15851,16277,15209,12945,8545,1665,3330,6660,13320,11347,7397,
                   14794,14295,11245,5017,10034,2599,5198,10396,5499,10998,4527,9054,767,1534,3068,
                   6136,12272,7075,14150,10959,4573,9146,823,1646,3292,6584,13168,8867,261,522,
                   1044,2088,4176,8352,1283,2566,5132,10264,5235,10470,5519,11038,4735,9470,3519,
                   7038,14076,10683,5941,11882,6295,12590,9759,2173,4346,8692,1963,3926,7852,15704,
                   16115,14757,14089,10833,4321,8642,1991,3982,7964,15928,14387,13349,11273,7249,14498,
                   13575,11853,6361,12722,10023,2573,5146,10292,5163,10326,5359,10718,6143,12286,7103,
                   14206,10943,4413,8826,183,366,732,1464,2928,5856,11712,8131,16262,15183,13021,
                   8697,1969,3938,7876,15752,16211,15077,12681,10065,2785,5570,11140,4939,9878,2415,
                   4830,9660,3899,7798,15596,15771,16245,15017,12561,9825,2177,4354,8708,75,150,
                   300,600,1200,2400,4800,9600,3907,7814,15628,15963,14581,13737,12049,6753,13506,
                   11719,8141,16282,15223,12973,8473,1649,3298,6596,13192,9043,741,1482,2964,5928,
                   11856,6371,12742,10191,3037,6074,12148,6827,13654,12015,6557,13114,8759,45,90,
                   180,360,720,1440,2880,5760,11520,7747,15494,15695,16093,14841,14257,11041,4609,
                   9218,3143,6286,12572,9851,2229,4458,8916,491,982,1964,3928,7856,15712,16003,
                   14661,14025,10705,6113,12226,7111,14222,11103,4861,9722,4023,8046,16092,14843,14261,
                   11049,4625,9250,3079,6158,12316,9339,3253,6506,13012,8683,1941,3882,7764,15528,
                   15635,15973,14473,13649,12001,6529,13058,8775,205,410,820,1640,3280,6560,13120,
                   8899,453,906,1812,3624,7248,14496,13571,11845,6345,12690,10087,2701,5402,10804,
                   4139,8278,1263,2526,5052,10104,2739,5478,10956,4571,9142,815,1630,3260,6520,
                   13040,8611,1797,3594,7188,14376,13331,11365,7305,14610,13927,10381,5465,10930,4391,
                   8782,223,446,892,1784,3568,7136,14272,11203,5061,10122,2903,5806,11612,7931,
                   15862,16303,15133,12921,8369,1313,2626,5252,10504,5715,11430,7439,14878,12415,9405,
                   3385,6770,13540,11659,8021,16042,14615,13933,10393,5489,10978,4487,8974,607,1214,
                   2428,4856,9712,4003,8006,16012,14683,14069,10665,5905,11810,6151,12302,9311,3325,
                   6650,13300,9131,789,1578,3156,6312,12624,9955,2437,4874,9748,2155,4310,8620,
                   1819,3638,7276,14552,13811,12197,6921,13842,10343,5261,10522,5751,11502,7583,15166,
                   12863,8253,1081,2162,4324,8648,2003,4006,8012,16024,14707,13989,10505,5713,11426,
                   7431,14862,12383,9469,3513,7026,14052,10635,5973,11946,6423,12846,8223,1149,2298,
                   4596,9192,915,1830,3660,7320,14640,13859,10245,5193,10386,5479,10958,4575,9150,
                   831,1662,3324,6648,13296,9123,773,1546,3092,6184,12368,9443,3461,6922,13844,
                   10347,5269,10538,5655,11310,7199,14398,13375,11325,7225,14450,13479,11533,7769,15538,
                   15655,15885,14425,13553,11681,7937,15874,14407,13517,11737,8177,16354,15239,13133,8921,
                   497,994,1988,3976,7952,15904,14339,13381,11465,7633,15266,13063,8781,217,434,
                   868,1736,3472,6944,13888,10435,5573,11146,4951,9902,2335,4670,9340,3259,6518,
                   13036,8603,1909,3818,7636,15272,13075,8805,137,274,548,1096,2192,4384,8768,
                   195,390,780,1560,3120,6240,12480,9667,4037,8074,16148,14955,12437,9577,3729,
                   7458,14916,12491,9685,4073,8146,16292,15115,12885,8425,1425,2850,5700,11400,7507,
                   15014,12559,9821,2297,4594,9188,907,1814,3628,7256,14512,13603,11781,6217,12434,
                   9575,3725,7450,14900,12331,9237,3177,6354,12708,9995,2645,5290,10580,5867,11734,
                   8175,16350,15359,13245,9017,561,1122,2244,4488,8976,611,1222,2444,4888,9776,
                   2083,4166,8332,1371,2742,5484,10968,4595,9190,911,1822,3644,7288,14576,13731,
                   12037,6729,13458,11623,7821,15642,15991,14509,13593,11889,6305,12610,9927,2509,5018,
                   10036,2603,5206,10412,5403,10806,4143,8286,1279,2558,5116,10232,2995,5990,11980,
                   6619,13238,9007,541,1082,2164,4328,8656,2019,4038,8076,16152,14963,12453,9481,
                   3665,7330,14660,14027,10709,6121,12242,7143,14286,11231,5117,10234,2999,5998,11996,
                   6651,13302,9135,797,1594,3188,6376,12752,10211,2949,5898,11796,6251,12502,9711,
                   3997,7994,15988,14507,13589,11881,6289,12578,9735,2125,4250,8500,1579,3158,6316,
                   12632,9971,2469,4938,9876,2411,4822,9644,3867,7734,15468,15515,15733,16041,14609,
                   13921,10369,5441,10882,4423,8846,351,702,1404,2808,5616,11232,4995,9990,2639,
                   5278,10556,5691,11382,7343,14686,14079,10685,5945,11890,6311,12622,9951,2557,5114,
                   10228,2987,5974,11948,6427,12854,8239,1053,2106,4212,8424,1427,2854,5708,11416,
                   7539,15078,12687,10077,2809,5618,11236,5003,10006,2671,5342,10684,5947,11894,6319,
                   12638,9983,2493,4986,9972,2475,4950,9900,2331,4662,9324,3227,6454,12908,8347,
                   1397,2794,5588,11176,4883,9766,2063,4126,8252,1083,2166,4332,8664,2035,4070,
                   8140,16280,15219,12965,8457,1617,3234,6468,12936,8531,1765,3530,7060,14120,10771,
                   4197,8394,1495,2990,5980,11960,6451,12902,8335,1373,2746,5492,10984,4499,8998,
                   527,1054,2108,4216,8432,1443,2886,5772,11544,7795,15590,15759,16221,15097,12721,
                   10017,2561,5122,10244,5195,10390,5487,10974,4607,9214,959,1918,3836,7672,15344,
                   13219,8965,585,1170,2340,4680,9360,3427,6854,13708,12123,6901,13802,12183,7021,
                   14042,10743,6061,12122,6903,13806,12191,7037,14074,10679,5933,11866,6391,12782,10143,
                   2941,5882,11764,8107,16214,15087,12701,10105,2737,5474,10948,4555,9110,879,1758,
                   3516,7032,14064,10659,5893,11786,6231,12462,9503,3709,7418,14836,14251,11029,4713,
                   9426,3559,7118,14236,11131,4789,9578,3735,7470,14940,12539,9653,3881,7762,15524,
                   15627,15957,14569,13713,12129,6785,13570,11847,6349,12698,10103,2733,5466,10932,4395,
                   8790,239,478,956,1912,3824,7648,15296,13251,9157,969,1938,3876,7752,15504,
                   15715,16005,14665,14033,10721,6017,12034,6727,13454,11615,7933,15866,16311,15149,12825,
                   8305,1185,2370,4740,9480,3667,7334,14668,14043,10741,6057,12114,6887,13774,12255,
                   7165,14330,11191,4909,9818,2295,4590,9180,1019,2038,4076,8152,16304,15139,12805,
                   8265,1233,2466,4932,9864,2387,4774,9548,3803,7606,15212,12955,8565,1705,3410,
                   6820,13640,11987,6629,13258,9175,1005,2010,4020,8040,16080,14819,14213,11081,4817,
                   9634,3847,7694,15388,15483,15541,15657,15889,14433,13441,11585,7873,15746,16199,15053,
                   12761,10225,2977,5954,11908,6475,12950,8559,1693,3386,6772,13544,11667,8037,16074,
                   14807,14317,11161,4977,9954,2439,4878,9756,2171,4342,8684,1947,3894,7788,15576,
                   15859,16293,15113,12881,8417,1409,2818,5636,11272,7251,14502,13583,11869,6393,12786,
                   10151,2829,5658,11316,7211,14422,13551,11677,8057,16114,14759,14093,10841,4337,8674,
                   1927,3854,7708,15416,15411,15397,15369,15441,15585,15745,16193,15041,12737,10177,3009,
                   6018,12036,6731,13462,11631,7837,15674,15927,14381,13337,11377,7329,14658,14023,10701,
                   6105,12210,6951,13902,10463,5629,11258,5047,10094,2719,5438,10876,4283,8566,1711,
                   3422,6844,13688,11955,6437,12874,8407,1517,3034,6068,12136,6803,13606,11791,6237,
                   12474,9527,3629,7258,14516,13611,11797,6249,12498,9703,3981,7962,15924,14379,13333,
                   11369,7313,14626,13831,10317,5337,10674,5927,11854,6367,12734,10047,2621,5242,10484,
                   5547,11094,4847,9694,4095,8190,16380,15291,13109,8745,17,34,68,136,272,
                   544,1088,2176,4352,8704,67,134,268,536,1072,2144,4288,8576,1859,3718,
                   7436,14872,12403,9381,3337,6674,13348,11275,7253,14506,13591,11885,6297,12594,9767,
                   2061,4122,8244,1067,2134,4268,8536,1779,3558,7116,14232,11123,4773,9546,3799,
                   7598,15196,13051,8629,1833,3666,7332,14664,14035,10725,6025,12050,6759,13518,11743,
                   8189,16378,15287,13101,8729,113,226,452,904,1808,3616,7232,14464,13635,11973,
                   6601,13202,9063,653,1306,2612,5224,10448,5603,11206,5071,10142,2943,5886,11772,
                   8123,16246,15023,12573,9849,2225,4450,8900,459,918,1836,3672,7344,14688,13955,
                   10565,5833,11666,8039,16078,14815,14333,11193,4913,9826,2183,4366,8732,123,246,
                   492,984,1968,3936,7872,15744,16195,15045,12745,10193,3041,6082,12164,6987,13974,
                   10607,5789,11578,7735,15470,15519,15741,16057,14641,13857,10241,5185,10370,5447,10894,
                   4447,8894,319,638,1276,2552,5104,10208,2947,5894,11788,6235,12470,9519,3613,
                   7226,14452,13483,11541,7785,15570,15847,16269,15193,13041,8609,1793,3586,7172,14344,
                   13395,11493,7561,15122,12903,8333,1369,2738,5476,10952,4563,9126,783,1566,3132,
                   6264,12528,9635,3845,7690,15380,15467,15509,15721,16017,14689,13953,10561,5825,11650,
                   8007,16014,14687,14077,10681,5937,11874,6279,12558,9823,2301,4602,9204,939,1878,
                   3756,7512,15024,12579,9733,2121,4242,8484,1547,3094,6188,12376,9459,3493,6986,
                   13972,10603,5781,11562,7703,15406,15391,15485,15545,15665,15905,14337,13377,11457,7617,
                   15234,13127,8909,473,946,1892,3784,7568,15136,12803,8261,1225,2450,4900,9800,
                   2259,4518,9036,731,1462,2924,5848,11696,7971,15942,14543,13789,12281,7089,14178,
                   10887,4429,8858,375,750,1500,3000,6000,12000,6531,13062,8783,221,442,884,
                   1768,3536,7072,14144,10947,4549,9098,855,1710,3420,6840,13680,11939,6405,12810,
                   8279,1261,2522,5044,10088,2707,5414,10828,4315,8630,1839,3678,7356,14712,14003,
                   10533,5641,11282,7271,14542,13791,12285,7097,14194,10919,4365,8730,119,238,476,
                   952,1904,3808,7616,15232,13123,8901,457,914,1828,3656,7312,14624,13827,10309,
                   5321,10642,5991,11982,6623,13246,9023,573,1146,2292,4584,9168,995,1990,3980,
                   7960,15920,14371,13317,11337,7377,14754,14087,10829,4313,8626,1831,3662,7324,14648,
                   13875,10277,5129,10258,5223,10446,5599,11198,4927,9854,2239,4478,8956,443,886,
                   1772,3544,7088,14176,10883,4421,8842,343,686,1372,2744,5488,10976,4483,8966,
                   591,1182,2364,4728,9456,3491,6982,13964,10587,5877,11754,8087,16174,14879,12413,
                   9401,3377,6754,13508,11723,8149,16298,15127,12909,8345,1393,2786,5572,11144,4947,
                   9894,2319,4638,9276,3131,6262,12524,9627,3957,7914,15828,16363,15253,13161,8849,
                   353,706,1412,2824,5648,11296,7171,14342,13391,11485,7673,15346,13223,8973,601,
                   1202,2404,4808,9616,3939,7878,15756,16219,15093,12713,10001,2657,5314,10628,5963,
                   11926,6511,13022,8703,1981,3962,7924,15848,16275,15205,12937,8529,1761,3522,7044,
                   14088,10835,4325,8650,2007,4014,8028,16056,14643,13861,10249,5201,10402,5383,10766,
                   4191,8382,1343,2686,5372,10744,6067,12134,6799,13598,11903,6333,12666,9911,2349,
                   4698,9396,3371,6742,13484,11547,7797,15594,15767,16237,15001,12657,9889,2305,4610,
                   9220,3147,6294,12588,9755,2165,4330,8660,2027,4054,8108,16216,15091,12709,9993,
                   2641,5282,10564,5835,11670,8047,16094,14847,14269,11065,4657,9314,3207,6414,12828,
                   8315,1205,2410,4820,9640,3859,7718,15436,15579,15861,16297,15121,12897,8321,1345,
                   2690,5380,10760,4179,8358,1295,2590,5180,10360,5299,10598,5775,11550,7807,15614,
                   15807,16189,14905,12337,9249,3073,6146,12292,9291,3285,6570,13140,8939,405,810,
                   1620,3240,6480,12960,8451,1605,3210,6420,12840,8211,1125,2250,4500,9000,531,
                   1062,2124,4248,8496,1571,3142,6284,12568,9843,2213,4426,8852,363,726,1452,
                   2904,5808,11616,7811,15622,15951,14557,13817,12209,6945,13890,10439,5581,11162,4983,
                   9966,2463,4926,9852,2235,4470,8940,411,822,1644,3288,6576,13152,8835,325,
                   650,1300,2600,5200,10400,5379,10758,4175,8350,1407,2814,5628,11256,5043,10086,
                   2703,5406,10812,4155,8310,1199,2398,4796,9592,3763,7526,15052,12763,10229,2985,
                   5970,11940,6411,12822,8303,1181,2362,4724,9448,3475,6950,13900,10459,5621,11242,
                   5015,10030,2591,5182,10364,5307,10614,5807,11614,7935,15870,16319,15165,12857,8241,
                   1057,2114,4228,8456,1619,3238,6476,12952,8563,1701,3402,6804,13608,11795,6245,
                   12490,9687,4077,8154,16308,15147,12821,8297,1169,2338,4676,9352,3411,6822,13644,
                   11995,6645,13290,9111,877,1754,3508,7016,14032,10723,6021,12042,6743,13486,11551,
                   7805,15610,15799,16173,14873,12401,9377,3329,6658,13316,11339,7381,14762,14103,10861,
                   4249,8498,1575,3150,6300,12600,9779,2085,4170,8340,1387,2774,5548,11096,4851,
                   9702,3983,7966,15932,14395,13365,11305,7185,14370,13319,11341,7385,14770,14119,10765,
                   4185,8370,1319,2638,5276,10552,5683,11366,7311,14622,13951,10429,5433,10866,4263,
                   8526,1759,3518,7036,14072,10675,5925,11850,6359,12718,10015,2685,5370,10740,6059,
                   12118,6895,13790,12287,7101,14202,10935,4397,8794,247,494,988,1976,3952,7904,
                   15808,16323,15301,13257,9169,993,1986,3972,7944,15888,14435,13445,11593,7889,15778,
                   16135,14925,12505,9713,4001,8002,16004,14667,14037,10729,6033,12066,6663,13326,11359,
                   7421,14842,14263,11053,4633,9266,3111,6222,12444,9595,3765,7530,15060,12779,10133,
                   2921,5842,11684,7947,15894,14447,13469,11641,7857,15714,16007,14669,14041,10737,6049,
                   12098,6855,13710,12127,6909,13818,12215,6957,13914,10487,5549,11098,4855,9710,3999,
                   7998,15996,14523,13621,11817,6161,12322,9223,3149,6298,12596,9771,2069,4138,8276,
                   1259,2518,5036,10072,2803,5606,11212,5083,10166,2863,5726,11452,7483,14966,12463,
                   9501,3705,7410,14820,14219,11093,4841,9682,4071,8142,16284,15227,12981,8489,1553,
                   3106,6212,12424,9555,3813,7626,15252,13163,8853,361,722,1444,2888,5776,11552,
                   7683,15366,15439,15581,15865,16305,15137,12801,8257,1217,2434,4868,9736,2131,4262,
                   8524,1755,3510,7020,14040,10739,6053,12106,6871,13742,12063,6781,13562,11703,7981,
                   15962,14583,13741,12057,6769,13538,11655,8013,16026,14711,13997,10521,5745,11490,7559,
                   15118,12895,8445,1465,2930,5860,11720,8147,16294,15119,12893,8441,1457,2914,5828,
                   11656,8019,16038,14607,13917,10489,5553,11106,4743,9486,3679,7358,14716,14011,10549,
                   5673,11346,7399,14798,14303,11261,5049,10098,2727,5454,10908,4475,8950,431,862,
                   1724,3448,6896,13792,12163,6981,13962,10583,5869,11738,8183,16366,15263,13181,8889,
                   305,610,1220,2440,4880,9760,2051,4102,8204,1115,2230,4460,8920,499,998,
                   1996,3992,7984,15968,14467,13637,11977,6609,13218,8967,589,1178,2356,4712,9424,
                   3555,7110,14220,11099,4853,9706,3991,7982,15964,14587,13749,12073,6673,13346,11271,
                   7245,14490,13687,11949,6425,12850,8231,1037,2074,4148,8296,1171,2342,4684,9368,
                   3443,6886,13772,12251,7157,14314,11159,4973,9946,2551,5102,10204,3067,6134,12268,
                   7067,14134,10799,4125,8250,1079,2158,4316,8632,1843,3686,7372,14744,14195,10917,
                   4361,8722,103,206,412,824,1648,3296,6592,13184,9027,709,1418,2836,5672,
                   11344,7395,14790,14287,11229,5113,10226,2983,5966,11932,6523,13046,8623,1821,3642,
                   7284,14568,13715,12133,6793,13586,11879,6285,12570,9847,2221,4442,8884,299,598,
                   1196,2392,4784,9568,3715,7430,14860,12379,9461,3497,6994,13988,10507,5717,11434,
                   7447,14894,12319,9341,3257,6514,13028,8587,1877,3754,7508,15016,12563,9829,2185,
                   4370,8740,11,22,44,88,176,352,704,1408,2816,5632,11264,7235,14470,
                   13647,11997,6649,13298,9127,781,1562,3124,6248,12496,9699,3973,7946,15892,14443,
                   13461,11625,7825,15650,15879,14413,13529,11761,8097,16194,15047,12749,10201,3057,6114,
                   12228,7115,14230,11119,4765,9530,3639,7278,14556,13819,12213,6953,13906,10471,5517,
                   11034,4727,9454,3487,6974,13948,10427,5429,10858,4247,8494,1567,3134,6268,12536,
                   9651,3877,7754,15508,15723,16021,14697,13969,10593,5761,11522,7751,15502,15711,16125,
                   14777,14129,10785,4097,8194,1095,2190,4380,8760,51,102,204,408,816,1632,
                   3264,6528,13056,8771,197,394,788,1576,3152,6304,12608,9923,2501,5002,10004,
                   2667,5334,10668,5915,11830,6191,12382,9471,3517,7034,14068,10667,5909,11818,6167,
                   12334,9247,3197,6394,12788,10155,2837,5674,11348,7403,14806,14319,11165,4985,9970,
                   2471,4942,9884,2427,4854,9708,3995,7990,15980,14491,13685,11945,6417,12834,8199,
                   1101,2202,4404,8808,147,294,588,1176,2352,4704,9408,3523,7046,14092,10843,
                   4341,8682,1943,3886,7772,15544,15667,15909,14345,13393,11489,7553,15106,12871,8397,
                   1497,2994,5988,11976,6611,13222,8975,605,1210,2420,4840,9680,4067,8134,16268,
                   15195,13045,8617,1809,3618,7236,14472,13651,12005,6537,13074,8807,141,282,564,
                   1128,2256,4512,9024,707,1414,2828,5656,11312,7203,14406,13519,11741,8185,16370,
                   15271,13069,8793,241,482,964,1928,3856,7712,15424,15555,15813,16329,15313,13281,
                   9089,833,1666,3332,6664,13328,11363,7301,14602,13911,10477,5529,11058,4647,9294,
                   3295,6590,13180,8891,309,618,1236,2472,4944,9888,2307,4614,9228,3163,6326,
                   12652,9883,2421,4842,9684,4075,8150,16300,15131,12917,8361,1297,2594,5188,10376,
                   5459,10918,4367,8734,127,254,508,1016,2032,4064,8128,16256,15171,12997,8649,
                   2001,4002,8004,16008,14675,14053,10633,5969,11938,6407,12814,8287,1277,2554,5108,
                   10216,2963,5926,11852,6363,12726,10031,2589,5178,10356,5291,10582,5871,11742,8191,
                   16382,15295,13117,8761,49,98,196,392,784,1568,3136,6272,12544,9795,2245,
                   4490,8980,619,1238,2476,4952,9904,2339,4678,9356,3419,6838,13676,11931,6517,
                   13034,8599,1901,3802,7604,15208,12947,8549,1673,3346,6692,13384,11475,7653,15306,
                   13271,9197,921,1842,3684,7368,14736,14179,10885,4425,8850,359,718,1436,2872,
                   5744,11488,7555,15110,12879,8413,1529,3058,6116,12232,7123,14246,11023,4701,9402,
                   3383,6766,13532,11771,8117,16234,14999,12653,9881,2417,4834,9668,4043,8086,16172,
                   14875,12405,9385,3345,6690,13380,11467,7637,15274,13079,8813,153,306,612,1224,
                   2448,4896,9792,2243,4486,8972,603,1206,2412,4824,9648,3875,7750,15500,15707,
                   16117,14761,14097,10849,4225,8450,1607,3214,6428,12856,8243,1061,2122,4244,8488,
                   1555,3110,6220,12440,9587,3749,7498,14996,12651,9877,2409,4818,9636,3851,7702,
                   15404,15387,15477,15529,15633,15969,14465,13633,11969,6593,13186,9031,717,1434,2868,
                   5736,11472,7651,15302,13263,9181,1017,2034,4068,8136,16272,15203,12933,8521,1745,
                   3490,6980,13960,10579,5861,11722,8151,16302,15135,12925,8377,1329,2658,5316,10632,
                   5971,11942,6415,12830,8319,1213,2426,4852,9704,3987,7974,15948,14555,13813,12201,
                   6929,13858,10247,5197,10394,5495,10990,4511,9022,575,1150,2300,4600,9200,931,
                   1862,3724,7448,14896,12323,9221,3145,6290,12580,9739,2133,4266,8532,1771,3542,
                   7084,14168,10995,4517,9034,727,1454,2908,5816,11632,7843,15686,16079,14813,14329,
                   11185,4897,9794,2247,4494,8988,635,1270,2540,5080,10160,2851,5702,11404,7515,
                   15030,12591,9757,2169,4338,8676,1931,3862,7724,15448,15603,15781,16137,14929,12513,
                   9601,3905,7810,15620,15947,14549,13801,12177,7009,14018,10695,6093,12186,7031,14062,
                   10655,6013,12026,6583,13166,8863,381,762,1524,3048,6096,12192,6915,13830,10319,
                   5341,10682,5943,11886,6303,12606,9791,2109,4218,8436,1451,2902,5804,11608,7923,
                   15846,16271,15197,13049,8625,1825,3650,7300,14600,13907,10469,5513,11026,4711,9422,
                   3551,7102,14204,10939,4405,8810,151,302,604,1208,2416,4832,9664,4035,8070,
                   16140,14939,12533,9641,3857,7714,15428,15563,15829,16361,15249,13153,8833,321,642,
                   1284,2568,5136,10272,5123,10246,5199,10398,5503,11006,4543,9086,703,1406,2812,
                   5624,11248,5027,10054,2767,5534,11068,4667,9334,3247,6494,12988,8507,1589,3178,
                   6356,12712,10003,2661,5322,10644,5995,11990,6639,13278,9215,957,1914,3828,7656,
                   15312,13283,9093,841,1682,3364,6728,13456,11619,7813,15626,15959,14573,13721,12145,
                   6817,13634,11975,6605,13210,9079,685,1370,2740,5480,10960,4579,9158,975,1950,
                   3900,7800,15600,15779,16133,14921,12497,9697,3969,7938,15876,14411,13525,11753,8081,
                   16162,14855,12365,9433,3569,7138,14276,11211,5077,10154,2839,5678,11356,7419,14838,
                   14255,11037,4729,9458,3495,6990,13980,10619,5813,11626,7831,15662,15903,14461,13497,
                   11569,7713,15426,15559,15821,16345,15345,13217,8961,577,1154,2308,4616,9232,3171,
                   6342,12684,10075,2805,5610,11220,5099,10198,3055,6110,12220,6971,13942,10415,5405,
                   10810,4151,8302,1183,2366,4732,9464,3507,7014,14028,10715,6133,12266,7063,14126,
                   10783,4221,8442,1463,2926,5852,11704,7987,15974,14479,13661,12025,6577,13154,8839,
                   333,666,1332,2664,5328,10656,5891,11782,6223,12446,9599,3773,7546,15092,12715,
                   10005,2665,5330,10660,5899,11798,6255,12510,9727,4029,8058,16116,14763,14101,10857,
                   4241,8482,1543,3086,6172,12344,9267,3109,6218,12436,9579,3733,7466,14932,12523,
                   9621,3945,7890,15780,16139,14933,12521,9617,3937,7874,15748,16203,15061,12777,10129,
                   2913,5826,11652,8011,16022,14703,13981,10617,5809,11618,7815,15630,15967,14589,13753,
                   12081,6689,13378,11463,7629,15258,13175,8877,281,562,1124,2248,4496,8992,515,
                   1030,2060,4120,8240,1059,2118,4236,8472,1651,3302,6604,13208,9075,677,1354,
                   2708,5416,10832,4323,8646,1999,3998,7996,15992,14515,13605,11785,6225,12450,9479,
                   3661,7322,14644,13867,10261,5225,10450,5607,11214,5087,10174,2879,5758,11516,7611,
                   15222,12975,8477,1657,3314,6628,13256,9171,997,1994,3988,7976,15952,14563,13701,
                   12105,6865,13730,12039,6733,13466,11639,7853,15706,16119,14765,14105,10865,4257,8514,
                   1735,3470,6940,13880,10291,5157,10314,5335,10670,5919,11838,6207,12414,9407,3389,
                   6778,13556,11691,7957,15914,14359,13421,11417,7537,15074,12679,10061,2777,5554,11108,
                   4747,9494,3695,7390,14780,14139,10805,4137,8274,1255,2510,5020,10040,2611,5222,
                   10444,5595,11190,4911,9822,2303,4606,9212,955,1910,3820,7640,15280,13091,8709,
                   73,146,292,584,1168,2336,4672,9344,3395,6790,13580,11867,6389,12778,10135,
                   2925,5850,11700,7979,15958,14575,13725,12153,6833,13666,11911,6477,12954,8567,1709,
                   3418,6836,13672,11923,6501,13002,8663,2029,4058,8116,16232,14995,12645,9865,2385,
                   4770,9540,3787,7574,15148,12827,8309,1193,2386,4772,9544,3795,7590,15180,13019,
                   8693,1961,3922,7844,15688,16083,14821,14217,11089,4833,9666,4039,8078,16156,14971,
                   12469,9513,3601,7202,14404,13515,11733,8169,16338,15335,13197,9049,753,1506,3012,
                   6024,12048,6755,13510,11727,8157,16314,15159,12845,8217,1137,2274,4548,9096,851,
                   1702,3404,6808,13616,11811,6149,12298,9303,3309,6618,13236,9003,533,1066,2132,
                   4264,8528,1763,3526,7052,14104,10867,4261,8522,1751,3502,7004,14008,10547,5669,
                   11338,7383,14766,14111,10877,4281,8562,1703,3406,6812,13624,11827,6181,12362,9431,
                   3565,7130,14260,11051,4629,9258,3095,6190,12380,9467,3509,7018,14036,10731,6037,
                   12074,6679,13358,11295,7293,14586,13751,12077,6681,13362,11303,7181,14362,13431,11437,
                   7449,14898,12327,9229,3161,6322,12644,9867,2389,4778,9556,3819,7638,15276,13083,
                   8821,169,338,676,1352,2704,5408,10816,4291,8582,1871,3742,7484,14968,12467,
                   9509,3593,7186,14372,13323,11349,7401,14802,14311,11149,4953,9906,2343,4686,9372,
                   3451,6902,13804,12187,7029,14058,10647,5997,11994,6647,13294,9119,893,1786,3572,
                   7144,14288,11235,4997,9994,2647,5294,10588,5883,11766,8111,16222,15103,12733,10041,
                   2609,5218,10436,5579,11158,4975,9950,2559,5118,10236,3003,6006,12012,6555,13110,
                   8751,29,58,116,232,464,928,1856,3712,7424,14848,12355,9413,3529,7058,
                   14116,10763,4181,8362,1303,2606,5212,10424,5427,10854,4239,8478,1663,3326,6652,
                   13304,9139,805,1610,3220,6440,12880,8419,1413,2826,5652,11304,7187,14374,13327,
                   11357,7417,14834,14247,11021,4697,9394,3367,6734,13468,11643,7861,15722,16023,14701,
                   13977,10609,5793,11586,7879,15758,16223,15101,12729,10033,2593,5186,10372,5451,10902,
                   4463,8926,511,1022,2044,4088,8176,16352,15235,13125,8905,465,930,1860,3720,
                   7440,14880,12291,9285,3273,6546,13092,8715,85,170,340,680,1360,2720,5440,
                   10880,4419,8838,335,670,1340,2680,5360,10720,6019,12038,6735,13470,11647,7869,
                   15738,16055,14637,13849,10353,5281,10562,5831,11662,8031,16062,14655,13885,10297,5169,
                   10338,5255,10510,5727,11454,7487,14974,12479,9533,3641,7282,14564,13707,12117,6889,
                   13778,12263,7053,14106,10871,4269,8538,1783,3566,7132,14264,11059,4645,9290,3287,
                   6574,13148,8955,437,874,1748,3496,6992,13984,10499,5701,11402,7511,15022,12575,
                   9853,2233,4466,8932,395,790,1580,3160,6320,12640,9859,2373,4746,9492,3691,
                   7382,14764,14107,10869,4265,8530,1767,3534,7068,14136,10803,4133,8266,1239,2478,
                   4956,9912,2355,4710,9420,3547,7094,14188,10907,4469,8938,407,814,1628,3256,
                   6512,13024,8579,1861,3722,7444,14888,12307,9317,3209,6418,12836,8203,1109,2218,
                   4436,8872,275,550,1100,2200,4400,8800,131,262,524,1048,2096,4192,8384,
                   1475,2950,5900,11800,6259,12518,9615,3933,7866,15732,16043,14613,13929,10385,5473,
                   10946,4551,9102,863,1726,3452,6904,13808,12195,6917,13834,10327,5357,10714,6135,
                   12270,7071,14142,10815,4157,8314,1207,2414,4828,9656,3891,7782,15564,15835,16373,
                   15273,13073,8801,129,258,516,1032,2064,4128,8256,1219,2438,4876,9752,2163,
                   4326,8652,2011,4022,8044,16088,14835,14245,11017,4689,9378,3335,6670,13340,11387,
                   7349,14698,13975,10605,5785,11570,7719,15438,15583,15869,16313,15153,12833,8193,1089,
                   2178,4356,8712,83,166,332,664,1328,2656,5312,10624,5955,11910,6479,12958,
                   8575,1725,3450,6900,13800,12179,7013,14026,10711,6125,12250,7159,14318,11167,4989,
                   9978,2487,4974,9948,2555,5110,10220,2971,5942,11884,6299,12598,9775,2077,4154,
                   8308,1195,2390,4780,9560,3827,7654,15308,13275,9205,937,1874,3748,7496,14992,
                   12643,9861,2377,4754,9508,3595,7190,14380,13339,11381,7337,14674,14055,10637,5977,
                   11954,6439,12878,8415,1533,3066,6132,12264,7059,14118,10767,4189,8378,1335,2670,
                   5340,10680,5939,11878,6287,12574,9855,2237,4474,8948,427,854,1708,3416,6832,
                   13664,11907,6469,12938,8535,1773,3546,7092,14184,10899,4453,8906,471,942,1884,
                   3768,7536,15072,12675,10053,2761,5522,11044,4619,9238,3183,6366,12732,10043,2613,
                   5226,10452,5611,11222,5103,10206,3071,6142,12284,7099,14198,10927,4381,8762,55,
                   110,220,440,880,1760,3520,7040,14080,10819,4293,8586,1879,3758,7516,15032,
                   12595,9765,2057,4114,8228,1035,2070,4140,8280,1267,2534,5068,10136,2931,5862,
                   11724,8155,16310,15151,12829,8313,1201,2402,4804,9608,3923,7846,15692,16091,14837,
                   14249,11025,4705,9410,3527,7054,14108,10875,4277,8554,1687,3374,6748,13496,11571,
                   7717,15434,15575,15853,16281,15217,12961,8449,1601,3202,6404,12808,8275,1253,2506,
                   5012,10024,2579,5158,10316,5339,10678,5935,11870,6399,12798,10175,2877,5754,11508,
                   7595,15190,13039,8605,1913,3826,7652,15304,13267,9189,905,1810,3620,7240,14480,
                   13667,11909,6473,12946,8551,1677,3354,6708,13416,11411,7525,15050,12759,10221,2969,
                   5938,11876,6283,12566,9839,2205,4410,8820,171,342,684,1368,2736,5472,10944,
                   4547,9094,847,1694,3388,6776,13552,11683,7941,15882,14423,13549,11673,8049,16098,
                   14727,14157,10969,4593,9186,903,1806,3612,7224,14448,13475,11525,7753,15506,15719,
                   16013,14681,14065,10657,5889,11778,6215,12430,9567,3837,7674,15348,13227,8981,617,
                   1234,2468,4936,9872,2403,4806,9612,3931,7862,15724,16027,14709,13993,10513,5729,
                   11458,7623,15246,13151,8957,441,882,1764,3528,7056,14112,10755,4165,8330,1367,
                   2734,5468,10936,4403,8806,143,286,572,1144,2288,4576,9152,963,1926,3852,
                   7704,15408,15395,15365,15433,15569,15841,16257,15169,12993,8641,1985,3970,7940,15880,
                   14419,13541,11657,8017,16034,14599,13901,10457,5617,11234,4999,9998,2655,5310,10620,
                   5819,11638,7855,15710,16127,14781,14137,10801,4129,8258,1223,2446,4892,9784,2099,
                   4198,8396,1499,2998,5996,11992,6643,13286,9103,861,1722,3444,6888,13776,12259,
                   7045,14090,10839,4333,8666,2039,4078,8156,16312,15155,12837,8201,1105,2210,4420,
                   8840,339,678,1356,2712,5424,10848,4227,8454,1615,3230,6460,12920,8371,1317,
                   2634,5268,10536,5651,11302,7183,14366,13439,11453,7481,14962,12455,9485,3673,7346,
                   14692,13963,10581,5865,11730,8167,16334,15327,13309,9145,817,1634,3268,6536,13072,
                   8803,133,266,532,1064,2128,4256,8512,1731,3462,6924,13848,10355,5285,10570,
                   5847,11694,7967,15934,14399,13373,11321,7217,14434,13447,11597,7897,15794,16167,14861,
                   12377,9457,3489,6978,13956,10571,5845,11690,7959,15918,14367,13437,11449,7473,14946,
                   12423,9549,3801,7602,15204,12939,8533,1769,3538,7076,14152,10963,4581,9162,983,
                   1966,3932,7864,15728,16035,14597,13897,10449,5601,11202,5063,10126,2911,5822,11644,
                   7867,15734,16047,14621,13945,10417,5409,10818,4295,8590,1887,3774,7548,15096,12723,
                   10021,2569,5138,10276,5131,10262,5231,10462,5631,11262,5055,10110,2751,5502,11004,
                   4539,9078,687,1374,2748,5496,10992,4515,9030,719,1438,2876,5752,11504,7587,
                   15174,13007,8669,2041,4082,8164,16328,15315,13285,9097,849,1698,3396,6792,13584,
                   11875,6277,12554,9815,2285,4570,9140,811,1622,3244,6488,12976,8483,1541,3082,
                   6164,12328,9235,3173,6346,12692,10091,2709,5418,10836,4331,8662,2031,4062,8124,
                   16248,15027,12581,9737,2129,4258,8516,1739,3478,6956,13912,10483,5541,11082,4823,
                   9646,3871,7742,15484,15547,15669,15913,14353,13409,11393,7489,14978,12615,9933,2521,
                   5042,10084,2699,5398,10796,4123,8246,1071,2142,4284,8568,1715,3430,6860,13720,
                   12147,6821,13642,11991,6637,13274,9207,941,1882,3764,7528,15056,12771,10117,2889,
                   5778,11556,7691,15382,15471,15517,15737,16049,14625,13825,10305,5313,10626,5959,11918,
                   6495,12990,8511,1597,3194,6388,12776,10131,2917,5834,11668,8043,16086,14831,14237,
                   11129,4785,9570,3719,7438,14876,12411,9397,3369,6738,13476,11531,7765,15530,15639,
                   15981,14489,13681,11937,6401,12802,8263,1229,2458,4916,9832,2195,4390,8780,219,
                   438,876,1752,3504,7008,14016,10691,6085,12170,6999,13998,10527,5757,11514,7607,
                   15214,12959,8573,1721,3442,6884,13768,12243,7141,14282,11223,5101,10202,3063,6126,
                   12252,7163,14326,11183,4893,9786,2103,4206,8412,1531,3062,6124,12248,7155,14310,
                   11151,4957,9914,2359,4718,9436,3579,7158,14316,11163,4981,9962,2455,4910,9820,
                   2299,4598,9196,923,1846,3692,7384,14768,14115,10757,4169,8338,1383,2766,5532,
                   11064,4659,9318,3215,6430,12860,8251,1077,2154,4308,8616,1811,3622,7244,14488,
                   13683,11941,6409,12818,8295,1165,2330,4660,9320,3219,6438,12876,8411,1525,3050,
                   6100,12200,6931,13862,10255,5213,10426,5431,10862,4255,8510,1599,3198,6396,12792,
                   10163,2853,5706,11412,7531,15062,12783,10141,2937,5874,11748,8075,16150,14959,12445,
                   9593,3761,7522,15044,12747,10197,3049,6098,12196,6923,13846,10351,5277,10554,5687,
                   11374,7327,14654,13887,10301,5177,10354,5287,10574,5855,11710,7999,15998,14527,13629,
                   11833,6193,12386,9351,3405,6810,13620,11819,6165,12330,9239,3181,6362,12724,10027,
                   2581,5162,10324,5355,10710,6127,12254,7167,14334,11199,4925,9850,2231,4462,8924,
                   507,1014,2028,4056,8112,16224,14979,12613,9929,2513,5026,10052,2763,5526,11052,
                   4635,9270,3119,6238,12476,9531,3637,7274,14548,13803,12181,7017,14034,10727,6029,
                   12058,6775,13550,11679,8061,16122,14775,14125,10777,4209,8418,1415,2830,5660,11320,
                   7219,14438,13455,11613,7929,15858,16295,15117,12889,8433,1441,2882,5764,11528,7763,
                   15526,15631,15965,14585,13745,12065,6657,13314,11335,7373,14746,14199,10925,4377,8754,
                   39,78,156,312,624,1248,2496,4992,9984,2627,5254,10508,5723,11446,7471,
                   14942,12543,9661,3897,7794,15588,15755,16213,15081,12689,10081,2689,5378,10756,4171,
                   8342,1391,2782,5564,11128,4787,9574,3727,7454,14908,12347,9269,3113,6226,12452,
                   9483,3669,7338,14676,14059,10645,5993,11986,6631,13262,9183,1021,2042,4084,8168,
                   16336,15331,13189,9033,721,1442,2884,5768,11536,7779,15558,15823,16349,15353,13233,
                   8993,513,1026,2052,4104,8208,1123,2246,4492,8984,627,1254,2508,5016,10032,
                   2595,5190,10380,5467,10934,4399,8798,255,510,1020,2040,4080,8160,16320,15299,
                   13253,9161,977,1954,3908,7816,15632,15971,14469,13641,11985,6625,13250,9159,973,
                   1946,3892,7784,15568,15843,16261,15177,13009,8673,1921,3842,7684,15368,15443,15589,
                   15753,16209,15073,12673,10049,2753,5506,11012,4683,9366,3439,6878,13756,12091,6709,
                   13418,11415,7533,15066,12791,10157,2841,5682,11364,7307,14614,13935,10397,5497,10994,
                   4519,9038,735,1470,2940,5880,11760,8099,16198,15055,12765,10233,2993,5986,11972,
                   6603,13206,9071,669,1338,2676,5352,10704,6115,12230,7119,14238,11135,4797,9594,
                   3767,7534,15068,12795,10165,2857,5714,11428,7435,14870,12399,9373,3449,6898,13796,
                   12171,6997,13994,10519,5741,11482,7671,15342,13215,9085,697,1394,2788,5576,11152,
                   4963,9926,2511,5022,10044,2619,5238,10476,5531,11062,4655,9310,3327,6654,13308,
                   9147,821,1642,3284,6568,13136,8931,389,778,1556,3112,6224,12448,9475,3653,
                   7306,14612,13931,10389,5481,10962,4583,9166,991,1982,3964,7928,15856,16291,15109,
                   12873,8401,1505,3010,6020,12040,6739,13478,11535,7773,15546,15671,15917,14361,13425,
                   11425,7425,14850,12359,9421,3545,7090,14180,10891,4437,8874,279,558,1116,2232,
                   4464,8928,387,774,1548,3096,6192,12384,9347,3397,6794,13588,11883,6293,12586,
                   9751,2157,4314,8628,1835,3670,7340,14680,14067,10661,5897,11794,6247,12494,9695,
                   4093,8186,16372,15275,13077,8809,145,290,580,1160,2320,4640,9280,3267,6534,
                   13068,8795,245,490,980,1960,3920,7840,15680,16067,14789,14281,11217,5089,10178,
                   3015,6030,12060,6779,13558,11695,7965,15930,14391,13357,11289,7281,14562,13703,12109,
                   6873,13746,12071,6669,13338,11383,7341,14682,14071,10669,5913,11826,6183,12366,9439,
                   3581,7162,14324,11179,4885,9770,2071,4142,8284,1275,2550,5100,10200,3059,6118,
                   12236,7131,14262,11055,4637,9274,3127,6254,12508,9723,4021,8042,16084,14827,14229,
                   11113,4753,9506,3591,7182,14364,13435,11445,7465,14930,12519,9613,3929,7858,15716,
                   16011,14677,14057,10641,5985,11970,6599,13198,9055,765,1530,3060,6120,12240,7139,
                   14278,11215,5085,10170,2871,5742,11484,7675,15350,13231,8989,633,1266,2532,5064,
                   10128,2915,5830,11660,8027,16054,14639,13853,10361,5297,10594,5767,11534,7775,15550,
                   15679,15933,14393,13361,11297,7169,14338,13383,11469,7641,15282,13095,8717,89,178,
                   356,712,1424,2848,5696,11392,7491,14982,12623,9949,2553,5106,10212,2955,5910,
                   11820,6171,12342,9263,3101,6202,12404,9387,3349,6698,13396,11499,7573,15146,12823,
                   8301,1177,2354,4708,9416,3539,7078,14156,10971,4597,9194,919,1838,3676,7352,
                   14704,13987,10501,5705,11410,7527,15054,12767,10237,3001,6002,12004,6539,13078,8815,
                   157,314,628,1256,2512,5024,10048,2755,5510,11020,4699,9398,3375,6750,13500,
                   11579,7733,15466,15511,15725,16025,14705,13985,10497,5697,11394,7495,14990,12639,9981,
                   2489,4978,9956,2443,4886,9772,2075,4150,8300,1179,2358,4716,9432,3571,7142,
                   14284,11227,5109,10218,2967,5934,11868,6395,12790,10159,2845,5690,11380,7339,14678,
                   14063,10653,6009,12018,6567,13134,8927,509,1018,2036,4072,8144,16288,15107,12869,
                   8393,1489,2978,5956,11912,6483,12966,8463,1629,3258,6516,13032,8595,1893,3786,
                   7572,15144,12819,8293,1161,2322,4644,9288,3283,6566,13132,8923,501,1002,2004,
                   4008,8016,16032,14595,13893,10441,5585,11170,4871,9742,2143,4286,8572,1723,3446,
                   6892,13784,12275,7077,14154,10967,4589,9178,1015,2030,4060,8120,16240,15011,12549,
                   9801,2257,4514,9028,715,1430,2860,5720,11440,7459,14918,12495,9693,4089,8178,
                   16356,15243,13141,8937,401,802,1604,3208,6416,12832,8195,1093,2186,4372,8744,
                   19,38,76,152,304,608,1216,2432,4864,9728,2115,4230,8460,1627,3254,
                   6508,13016,8691,1957,3914,7828,15656,15891,14437,13449,11601,7905,15810,16327,15309,
                   13273,9201,929,1858,3716,7432,14864,12387,9349,3401,6802,13604,11787,6229,12458,
                   9495,3693,7386,14772,14123,10773,4201,8402,1511,3022,6044,12088,6707,13414,11407,
                   7517,15034,12599,9773,2073,4146,8292,1163,2326,4652,9304,3315,6630,13260,9179,
                   1013,2026,4052,8104,16208,15075,12677,10057,2769,5538,11076,4811,9622,3951,7902,
                   15804,16187,14901,12329,9233,3169,6338,12676,10059,2773,5546,11092,4843,9686,4079,
                   8158,16316,15163,12853,8233,1041,2082,4164,8328,1363,2726,5452,10904,4467,8934,
                   399,798,1596,3192,6384,12768,10115,2885,5770,11540,7787,15574,15855,16285,15225,
                   12977,8481,1537,3074,6148,12296,9299,3301,6602,13204,9067,661,1322,2644,5288,
                   10576,5859,11718,8143,16286,15231,12989,8505,1585,3170,6340,12680,10067,2789,5578,
                   11156,4971,9942,2543,5086,10172,2875,5750,11500,7579,15158,12847,8221,1145,2290,
                   4580,9160,979,1958,3916,7832,15664,15907,14341,13385,11473,7649,15298,13255,9165,
                   985,1970,3940,7880,15760,16227,14981,12617,9937,2529,5058,10116,2891,5782,11564,
                   7707,15414,15407,15389,15481,15537,15649,15873,14401,13505,11713,8129,16258,15175,13005,
                   8665,2033,4066,8132,16264,15187,13029,8585,1873,3746,7492,14984,12627,9957,2441,
                   4882,9764,2059,4118,8236,1051,2102,4204,8408,1523,3046,6092,12184,7027,14054,
                   10639,5981,11962,6455,12910,8351,1405,2810,5620,11240,5011,10022,2575,5150,10300,
                   5179,10358,5295,10590,5887,11774,8127,16254,15039,12605,9785,2097,4194,8388,1483,
                   2966,5932,11864,6387,12774,10127,2909,5818,11636,7851,15702,16111,14749,14201,10929,
                   4385,8770,199,398,796,1592,3184,6368,12736,10179,3013,6026,12052,6763,13526,
                   11759,8093,16186,14903,12333,9241,3185,6370,12740,10187,3029,6058,12116,6891,13782,
                   12271,7069,14138,10807,4141,8282,1271,2542,5084,10168,2867,5734,11468,7643,15286,
                   13103,8733,121,242,484,968,1936,3872,7744,15488,15683,16069,14793,14289,11233,
                   4993,9986,2631,5262,10524,5755,11510,7599,15198,13055,8637,1849,3698,7396,14792,
                   14291,11237,5001,10002,2663,5326,10652,6011,12022,6575,13150,8959,445,890,1780,
                   3560,7120,14240,11011,4677,9354,3415,6830,13660,12027,6581,13162,8855,365,730,
                   1460,2920,5840,11680,7939,15878,14415,13533,11769,8113,16226,14983,12621,9945,2545,
                   5090,10180,3019,6038,12076,6683,13366,11311,7197,14394,13367,11309,7193,14386,13351,
                   11277,7257,14514,13607,11789,6233,12466,9511,3597,7194,14388,13355,11285,7273,14546,
                   13799,12173,7001,14002,10535,5645,11290,7287,14574,13727,12157,6841,13682,11943,6413,
                   12826,8311,1197,2394,4788,9576,3731,7462,14924,12507,9717,4009,8018,16036,14603,
                   13909,10473,5521,11042,4615,9230,3167,6334,12668,9915,2357,4714,9428,3563,7126,
                   14252,11035,4725,9450,3479,6958,13916,10491,5557,11114,4759,9518,3615,7230,14460,
                   13499,11573,7721,15442,15591,15757,16217,15089,12705,9985,2625,5250,10500,5707,11414,
                   7535,15070,12799,10173,2873,5746,11492,7563,15126,12911,8349,1401,2802,5604,11208,
                   5075,10150,2831,5662,11324,7227,14454,13487,11549,7801,15602,15783,16141,14937,12529,
                   9633,3841,7682,15364,15435,15573,15849,16273,15201,12929,8513,1729,3458,6916,13832,
                   10323,5349,10698,6103,12206,6943,13886,10303,5181,10362,5303,10606,5791,11582,7743,
                   15486,15551,15677,15929,14385,13345,11265,7233,14466,13639,11981,6617,13234,8999,525,
                   1050,2100,4200,8400,1507,3014,6028,12056,6771,13542,11663,8029,16058,14647,13869,
                   10265,5233,10466,5511,11022,4703,9406,3391,6782,13564,11707,7989,15978,14487,13677,
                   11929,6513,13026,8583,1869,3738,7476,14952,12435,9573,3721,7442,14884,12299,9301,
                   3305,6610,13220,8971,597,1194,2388,4776,9552,3811,7622,15244,13147,8949,425,
                   850,1700,3400,6800,13600,11779,6213,12426,9559,3821,7642,15284,13099,8725,105,
                   210,420,840,1680,3360,6720,13440,11587,7877,15754,16215,15085,12697,10097,2721,
                   5442,10884,4427,8854,367,734,1468,2936,5872,11744,8067,16134,14927,12509,9721,
                   4017,8034,16068,14795,14293,11241,5009,10018,2567,5134,10268,5243,10486,5551,11102,
                   4863,9726,4031,8062,16124,14779,14133,10793,4113,8226,1031,2062,4124,8248,1075,
                   2150,4300,8600,1907,3814,7628,15256,13171,8869,265,530,1060,2120,4240,8480,
                   1539,3078,6156,12312,9331,3237,6474,12948,8555,1685,3370,6740,13480,11539,7781,
                   15562,15831,16365,15257,13169,8865,257,514,1028,2056,4112,8224,1027,2054,4108,
                   8216,1139,2278,4556,9112,883,1766,3532,7064,14128,10787,4101,8202,1111,2222,
                   4444,8888,307,614,1228,2456,4912,9824,2179,4358,8716,91,182,364,728,
                   1456,2912,5824,11648,8003,16006,14671,14045,10745,6065,12130,6791,13582,11871,6397,
                   12794,10167,2861,5722,11444,7467,14934,12527,9629,3961,7922,15844,16267,15189,13033,
                   8593,1889,3778,7556,15112,12883,8421,1417,2834,5668,11336,7379,14758,14095,10845,
                   4345,8690,1959,3918,7836,15672,15923,14373,13321,11345,7393,14786,14279,11213,5081,
                   10162,2855,5710,11420,7547,15094,12719,10013,2681,5362,10724,6027,12054,6767,13534,
                   11775,8125,16250,15031,12589,9753,2161,4322,8644,1995,3990,7980,15960,14579,13733,
                   12041,6737,13474,11527,7757,15514,15735,16045,14617,13937,10401,5377,10754,4167,8334,
                   1375,2750,5500,11000,4531,9062,655,1310,2620,5240,10480,5539,11078,4815,9630,
                   3967,7934,15868,16315,15157,12841,8209,1121,2242,4484,8968,595,1190,2380,4760,
                   9520,3619,7238,14476,13659,12021,6569,13138,8935,397,794,1588,3176,6352,12704,
                   9987,2629,5258,10516,5739,11478,7663,15326,13311,9149,825,1650,3300,6600,13200,
                   9059,645,1290,2580,5160,10320,5347,10694,6095,12190,7039,14078,10687,5949,11898,
                   6327,12654,9887,2429,4858,9716,4011,8022,16044,14619,13941,10409,5393,10786,4103,
                   8206,1119,2238,4476,8952,435,870,1740,3480,6960,13920,10371,5445,10890,4439,
                   8878,287,574,1148,2296,4592,9184,899,1798,3596,7192,14384,13347,11269,7241,
                   14482,13671,11917,6489,12978,8487,1549,3098,6196,12392,9363,3429,6858,13716,12139,
                   6805,13610,11799,6253,12506,9719,4013,8026,16052,14635,13845,10345,5265,10530,5639,
                   11278,7263,14526,13631,11837,6201,12402,9383,3341,6682,13364,11307,7189,14378,13335,
                   11373,7321,14642,13863,10253,5209,10418,5415,10830,4319,8638,1855,3710,7420,14840,
                   14259,11045,4617,9234,3175,6350,12700,10107,2741,5482,10964,4587,9174,1007,2014,
                   4028,8056,16112,14755,14085,10825,4305,8610,1799,3598,7196,14392,13363,11301,7177,
                   14354,13415,11405,7513,15026,12583,9741,2137,4274,8548,1675,3350,6700,13400,11507,
                   7589,15178,13015,8685,1945,3890,7780,15560,15827,16357,15241,13137,8929,385,770,
                   1540,3080,6160,12320,9219,3141,6282,12564,9835,2197,4394,8788,235,470,940,
                   1880,3760,7520,15040,12739,10181,3017,6034,12068,6667,13334,11375,7325,14650,13879,
                   10285,5145,10290,5159,10318,5343,10686,5951,11902,6335,12670,9919,2365,4730,9460,
                   3499,6998,13996,10523,5749,11498,7575,15150,12831,8317,1209,2418,4836,9672,4051,
                   8102,16204,15067,12789,10153,2833,5666,11332,7371,14742,14191,10909,4473,8946,423,
                   846,1692,3384,6768,13536,11651,8005,16010,14679,14061,10649,6001,12002,6535,13070,
                   8799,253,506,1012,2024,4048,8096,16192,15043,12741,10185,3025,6050,12100,6859,
                   13718,12143,6813,13626,11831,6189,12378,9463,3501,7002,14004,10539,5653,11306,7191,
                   14382,13343,11389,7353,14706,13991,10509,5721,11442,7463,14926,12511,9725,4025,8050,
                   16100,14731,14165,10985,4497,8994,519,1038,2076,4152,8304,1187,2374,4748,9496,
                   3699,7398,14796,14299,11253,5033,10066,2791,5582,11164,4987,9974,2479,4958,9916,
                   2363,4726,9452,3483,6966,13932,10395,5493,10986,4503,9006,543,1086,2172,4344,
                   8688,1955,3910,7820,15640,15987,14501,13577,11857,6369,12738,10183,3021,6042,12084,
                   6699,13398,11503,7581,15162,12855,8237,1049,2098,4196,8392,1491,2982,5964,11928,
                   6515,13030,8591,1885,3770,7540,15080,12691,10085,2697,5394,10788,4107,8214,1135,
                   2270,4540,9080,691,1382,2764,5528,11056,4643,9286,3279,6558,13116,8763,53,
                   106,212,424,848,1696,3392,6784,13568,11843,6341,12682,10071,2797,5594,11188,
                   4907,9814,2287,4574,9148,827,1654,3308,6616,13232,8995,517,1034,2068,4136,
                   8272,1251,2502,5004,10008,2675,5350,10700,6107,12214,6959,13918,10495,5565,11130,
                   4791,9582,3743,7486,14972,12475,9525,3625,7250,14500,13579,11861,6377,12754,10215,
                   2957,5914,11828,6187,12374,9455,3485,6970,13940,10411,5397,10794,4119,8238,1055,
                   2110,4220,8440,1459,2918,5836,11672,8051,16102,14735,14173,11001,4529,9058,647,
                   1294,2588,5176,10352,5283,10566,5839,11678,8063,16126,14783,14141,10809,4145,8290,
                   1159,2318,4636,9272,3123,6246,12492,9691,4085,8170,16340,15339,13205,9065,657,
                   1314,2628,5256,10512,5731,11462,7631,15262,13183,8893,313,626,1252,2504,5008,
                   10016,2563,5126,10252,5211,10422,5423,10846,4351,8702,1983,3966,7932,15864,16307,
                   15141,12809,8273,1249,2498,4996,9992,2643,5286,10572,5851,11702,7983,15966,14591,
                   13757,12089,6705,13410,11399,7501,15002,12663,9901,2329,4658,9316,3211,6422,12844,
                   8219,1141,2282,4564,9128,787,1574,3148,6296,12592,9763,2053,4106,8212,1131,
                   2262,4524,9048,755,1510,3020,6040,12080,6691,13382,11471,7645,15290,13111,8749,
                   25,50,100,200,400,800,1600,3200,6400,12800,8259,1221,2442,4884,9768,
                   2067,4134,8268,1243,2486,4972,9944,2547,5094,10188,3035,6070,12140,6811,13622,
                   11823,6173,12346,9271,3117,6234,12468,9515,3605,7210,14420,13547,11669,8041,16082,
                   14823,14221,11097,4849,9698,3975,7950,15900,14459,13493,11561,7697,15394,15367,15437,
                   15577,15857,16289,15105,12865,8385,1473,2946,5892,11784,6227,12454,9487,3677,7354,
                   14708,13995,10517,5737,11474,7655,15310,13279,9213,953,1906,3812,7624,15248,13155,
                   8837,329,658,1316,2632,5264,10528,5635,11270,7247,14494,13695,11965,6457,12914,
                   8359,1293,2586,5172,10344,5267,10534,5647,11294,7295,14590,13759,12093,6713,13426,
                   11431,7437,14874,12407,9389,3353,6706,13412,11403,7509,15018,12567,9837,2201,4402,
                   8804,139,278,556,1112,2224,4448,8896,451,902,1804,3608,7216,14432,13443,
                   11589,7881,15762,16231,14989,12633,9969,2465,4930,9860,2379,4758,9516,3611,7222,
                   14444,13467,11637,7849,15698,16103,14733,14169,10993,4513,9026,711,1422,2844,5688,
                   11376,7331,14662,14031,10717,6137,12274,7079,14158,10975,4605,9210,951,1902,3804,
                   7608,15216,12963,8453,1609,3218,6436,12872,8403,1509,3018,6036,12072,6675,13350,
                   11279,7261,14522,13623,11821,6169,12338,9255,3085,6170,12340,9259,3093,6186,12372,
                   9451,3477,6954,13908,10475,5525,11050,4631,9262,3103,6206,12412,9403,3381,6762,
                   13524,11755,8085,16170,14871,12397,9369,3441,6882,13764,12235,7125,14250,11031,4717,
                   9434,3575,7150,14300,11259,5045,10090,2711,5422,10844,4347,8694,1967,3934,7868,
                   15736,16051,14629,13833,10321,5345,10690,6087,12174,7007,14014,10559,5693,11386,7351,
                   14702,13983,10621,5817,11634,7847,15694,16095,14845,14265,11057,4641,9282,3271,6542,
                   13084,8827,181,362,724,1448,2896,5792,11584,7875,15750,16207,15069,12793,10161,
                   2849,5698,11396,7499,14998,12655,9885,2425,4850,9700,3979,7958,15916,14363,13429,
                   11433,7441,14882,12295,9293,3289,6578,13156,8843,341,682,1364,2728,5456,10912,
                   4355,8710,79,158,316,632,1264,2528,5056,10112,2883,5766,11532,7771,15542,
                   15663,15901,14457,13489,11553,7681,15362,15431,15565,15833,16369,15265,13057,8769,193,
                   386,772,1544,3088,6176,12352,9411,3525,7050,14100,10859,4245,8490,1559,3118,
                   6236,12472,9523,3621,7242,14484,13675,11925,6505,13010,8679,1933,3866,7732,15464,
                   15507,15717,16009,14673,14049,10625,5953,11906,6471,12942,8543,1789,3578,7156,14312,
                   11155,4965,9930,2519,5038,10076,2811,5622,11244,5019,10038,2607,5214,10428,5435,
                   10870,4271,8542,1791,3582,7164,14328,11187,4901,9802,2263,4526,9052,763,1526,
                   3052,6104,12208,6947,13894,10447,5597,11194,4919,9838,2207,4414,8828,187,374,
                   748,1496,2992,5984,11968,6595,13190,9039,733,1466,2932,5864,11728,8163,16326,
                   15311,13277,9209,945,1890,3780,7560,15120,12899,8325,1353,2706,5412,10824,4307,
                   8614,1807,3614,7228,14456,13491,11557,7689,15378,15463,15501,15705,16113,14753,14081,
                   10817,4289,8578,1863,3726,7452,14904,12339,9253,3081,6162,12324,9227,3157,6314,
                   12628,9963,2453,4906,9812,2283,4566,9132,795,1590,3180,6360,12720,10019,2565,
                   5130,10260,5227,10454,5615,11230,5119,10238,3007,6014,12028,6587,13174,8879,285,
                   570,1140,2280,4560,9120,771,1542,3084,6168,12336,9251,3077,6154,12308,9323,
                   3221,6442,12884,8427,1429,2858,5716,11432,7443,14886,12303,9309,3321,6642,13284,
                   9099,853,1706,3412,6824,13648,12003,6533,13066,8791,237,474,948,1896,3792,
                   7584,15168,12995,8645,1993,3986,7972,15944,14547,13797,12169,6993,13986,10503,5709,
                   11418,7543,15086,12703,10109,2745,5490,10980,4491,8982,623,1246,2492,4984,9968,
                   2467,4934,9868,2395,4790,9580,3739,7478,14956,12443,9589,3753,7506,15012,12555,
                   9813,2281,4562,9124,779,1558,3116,6232,12464,9507,3589,7178,14356,13419,11413,
                   7529,15058,12775,10125,2905,5810,11620,7819,15638,15983,14493,13689,11953,6433,12866,
                   8391,1485,2970,5940,11880,6291,12582,9743,2141,4282,8564,1707,3414,6828,13656,
                   12019,6565,13130,8919,493,986,1972,3944,7888,15776,16131,14917,12489,9681,4065,
                   8130,16260,15179,13013,8681,1937,3874,7748,15496,15699,16101,14729,14161,10977,4481,
                   8962,583,1166,2332,4664,9328,3235,6470,12940,8539,1781,3562,7124,14248,11027,
                   4709,9418,3543,7086,14172,11003,4533,9066,663,1326,2652,5304,10608,5795,11590,
                   7887,15774,16255,15037,12601,9777,2081,4162,8324,1355,2710,5420,10840,4339,8678,
                   1935,3870,7740,15480,15539,15653,15881,14417,13537,11649,8001,16002,14663,14029,10713,
                   6129,12258,7047,14094,10847,4349,8698,1975,3950,7900,15800,16179,14885,12297,9297,
                   3297,6594,13188,9035,725,1450,2900,5800,11600,7907,15814,16335,15325,13305,9137,
                   801,1602,3204,6408,12816,8291,1157,2314,4628,9256,3091,6182,12364,9435,3573,
                   7146,14292,11243,5013,10026,2583,5166,10332,5371,10742,6063,12126,6911,13822,12223,
                   6973,13946,10423,5421,10842,4343,8686,1951,3902,7804,15608,15795,16165,14857,12369,
                   9441,3457,6914,13828,10315,5333,10666,5911,11822,6175,12350,9279,3133,6266,12532,
                   9643,3861,7722,15444,15595,15765,16233,14993,12641,9857,2369,4738,9476,3659,7318,
                   14636,13851,10357,5289,10578,5863,11726,8159,16318,15167,12861,8249,1073,2146,4292,
                   8584,1875,3750,7500,15000,12659,9893,2313,4626,9252,3083,6166,12332,9243,3189,
                   6378,12756,10219,2965,5930,11860,6379,12758,10223,2973,5946,11892,6315,12630,9967,
                   2461,4922,9844,2219,4438,8876,283,566,1132,2264,4528,9056,643,1286,2572,
                   5144,10288,5155,10310,5327,10654,6015,12030,6591,13182,8895,317,634,1268,2536,
                   5072,10144,2819,5638,11276,7259,14518,13615,11805,6265,12530,9639,3853,7706,15412,
                   15403,15381,15465,15505,15713,16001,14657,14017,10689,6081,12162,6983,13966,10591,5885,
                   11770,8119,16238,15007,12669,9913,2353,4706,9412,3531,7062,14124,10779,4213,8426,
                   1431,2862,5724,11448,7475,14950,12431,9565,3833,7666,15332,13195,9045,745,1490,
                   2980,5960,11920,6499,12998,8655,2013,4026,8052,16104,14739,14181,10889,4433,8866,
                   263,526,1052,2104,4208,8416,1411,2822,5644,11288,7283,14566,13711,12125,6905,
                   13810,12199,6925,13850,10359,5293,10586,5879,11758,8095,16190,14911,12349,9273,3121,
                   6242,12484,9675,4053,8106,16212,15083,12693,10089,2705,5410,10820,4299,8598,1903,
                   3806,7612,15224,12979,8485,1545,3090,6180,12360,9427,3557,7114,14228,11115,4757,
                   9514,3607,7214,14428,13563,11701,7977,15954,14567,13709,12121,6897,13794,12167,6989,
                   13978,10615,5805,11610,7927,15854,16287,15229,12985,8497,1569,3138,6276,12552,9811,
                   2277,4554,9108,875,1750,3500,7000,14000,10531,5637,11274,7255,14510,13599,11901,
                   6329,12658,9895,2317,4634,9268,3115,6230,12460,9499,3701,7402,14804,14315,11157,
                   4969,9938,2535,5070,10140,2939,5878,11756,8091,16182,14895,12317,9337,3249,6498,
                   12996,8651,2005,4010,8020,16040,14611,13925,10377,5457,10914,4359,8718,95,190,
                   380,760,1520,3040,6080,12160,6979,13958,10575,5853,11706,7991,15982,14495,13693,
                   11961,6449,12898,8327,1357,2714,5428,10856,4243,8486,1551,3102,6204,12408,9395,
                   3365,6730,13460,11627,7829,15658,15895,14445,13465,11633,7841,15682,16071,14797,14297,
                   11249,5025,10050,2759,5518,11036,4731,9462,3503,7006,14012,10555,5685,11370,7319,
                   14638,13855,10365,5305,10610,5799,11598,7903,15806,16191,14909,12345,9265,3105,6210,
                   12420,9547,3797,7594,15188,13035,8597,1897,3794,7588,15176,13011,8677,1929,3858,
                   7716,15432,15571,15845,16265,15185,13025,8577,1857,3714,7428,14856,12371,9445,3465,
                   6930,13860,10251,5205,10410,5399,10798,4127,8254,1087,2174,4348,8696,1971,3942,
                   7884,15768,16243,15013,12553,9809,2273,4546,9092,843,1686,3372,6744,13488,11555,
                   7685,15370,15447,15597,15769,16241,15009,12545,9793,2241,4482,8964,587,1174,2348,
                   4696,9392,3363,6726,13452,11611,7925,15850,16279,15213,12953,8561,1697,3394,6788,
                   13576,11859,6373,12746,10199,3053,6106,12212,6955,13910,10479,5533,11066,4663,9326,
                   3231,6462,12924,8379,1333,2666,5332,10664,5907,11814,6159,12318,9343,3261,6522,
                   13044,8619,1813,3626,7252,14504,13587,11877,6281,12562,9831,2189,4378,8756,43,
                   86,172,344,688,1376,2752,5504,11008,4675,9350,3407,6814,13628,11835,6197,
                   12394,9367,3437,6874,13748,12075,6677,13354,11287,7277,14554,13815,12205,6937,13874,
                   10279,5133,10266,5239,10478,5535,11070,4671,9342,3263,6526,13052,8635,1845,3690,
                   7380,14760,14099,10853,4233,8466,1639,3278,6556,13112,8755,37,74,148,296,
                   592,1184,2368,4736,9472,3651,7302,14604,13915,10485,5545,11090,4839,9678,4063,
                   8126,16252,15035,12597,9769,2065,4130,8260,1227,2454,4908,9816,2291,4582,9164,
                   987,1974,3948,7896,15792,16163,14853,12361,9425,3553,7106,14212,11083,4821,9642,
                   3863,7726,15452,15611,15797,16169,14865,12385,9345,3393,6786,13572,11851,6357,12714,
                   10007,2669,5338,10676,5931,11862,6383,12766,10239,3005,6010,12020,6571,13142,8943,
                   413,826,1652,3304,6608,13216,8963,581,1162,2324,4648,9296,3299,6598,13196,
                   9051,757,1514,3028,6056,12112,6883,13766,12239,7133,14266,11063,4653,9306,3319,
                   6638,13276,9211,949,1898,3796,7592,15184,13027,8581,1865,3730,7460,14920,12499,
                   9701,3977,7954,15908,14347,13397,11497,7569,15138,12807,8269,1241,2482,4964,9928,
                   2515,5030,10060,2779,5558,11116,4763,9526,3631,7262,14524,13627,11829,6185,12370,
                   9447,3469,6938,13876,10283,5141,10282,5143,10286,5151,10302,5183,10366,5311,10622,
                   5823,11646,7871,15742,16063,14653,13881,10289,5153,10306,5319,10638,5983,11966,6463,
                   12926,8383,1341,2682,5364,10728,6035,12070,6671,13342,11391,7357,14714,14007,10541,
                   5657,11314,7207,14414,13535,11773,8121,16242,15015,12557,9817,2289,4578,9156,971,
                   1942,3884,7768,15536,15651,15877,14409,13521,11745,8065,16130,14919,12493,9689,4081,
                   8162,16324,15307,13269,9193,913,1826,3652,7304,14608,13923,10373,5449,10898,4455,
                   8910,479,958,1916,3832,7664,15328,13187,9029,713,1426,2852,5704,11408,7523,
                   15046,12751,10205,3065,6130,12260,7051,14102,10863,4253,8506,1591,3182,6364,12728,
                   10035,2597,5194,10388,5483,10966,4591,9182,1023,2046,4092,8184,16368,15267,13061,
                   8777,209,418,836,1672,3344,6688,13376,11459,7621,15242,13143,8941,409,818,
                   1636,3272,6544,13088,8707,69,138,276,552,1104,2208,4416,8832,323,646,
                   1292,2584,5168,10336,5251,10502,5711,11422,7551,15102,12735,10045,2617,5234,10468,
                   5515,11030,4719,9438,3583,7166,14332,11195,4917,9834,2199,4398,8796,251,502,
                   1004,2008,4016,8032,16064,14787,14277,11209,5073,10146,2823,5646,11292,7291,14582,
                   13743,12061,6777,13554,11687,7949,15898,14455,13485,11545,7793,15586,15751,16205,15065,
                   12785,10145,2817,5634,11268,7243,14486,13679,11933,6521,13042,8615,1805,3610,7220,
                   14440,13459,11621,7817,15634,15975,14477,13657,12017,6561,13122,8903,461,922,1844,
                   3688,7376,14752,14083,10821,4297,8594,1895,3790,7580,15160,12851,8229,1033,2066,
                   4132,8264,1235,2470,4940,9880,2419,4838,9676,4059,8118,16236,15003,12661,9897,
                   2321,4642,9284,3275,6550,13100,8731,117,234,468,936,1872,3744,7488,14976,
                   12611,9925,2505,5010,10020,2571,5142,10284,5147,10294,5167,10334,5375,10750,6079,
                   12158,6847,13694,11967,6461,12922,8375,1325,2650,5300,10600,5779,11558,7695,15390,
                   15487,15549,15673,15921,14369,13313,11329,7361,14722,14151,10957,4569,9138,807,1614,
                   3228,6456,12912,8355,1285,2570,5140,10280,5139,10278,5135,10270,5247,10494,5567,
                   11134,4799,9598,3775,7550,15100,12731,10037,2601,5202,10404,5387,10774,4207,8414,
                   1535,3070,6140,12280,7091,14182,10895,4445,8890,311,622,1244,2488,4976,9952,
                   2435,4870,9740,2139,4278,8556,1691,3382,6764,13528,11763,8101,16202,15063,12781,
                   10137,2929,5858,11716,8139,16278,15215,12957,8569,1713,3426,6852,13704,12115,6885,
                   13770,12247,7149,14298,11255,5037,10074,2807,5614,11228,5115,10230,2991,5982,11964,
                   6459,12918,8367,1309,2618,5236,10472,5523,11046,4623,9246,3199,6398,12796,10171,
                   2869,5738,11476,7659,15318,13295,9117,889,1778,3556,7112,14224,11107,4741,9482,
                   3671,7342,14684,14075,10677,5929,11858,6375,12750,10207,3069,6138,12276,7083,14166,
                   10991,4509,9018,567,1134,2268,4536,9072,675,1350,2700,5400,10800,4131,8262,
                   1231,2462,4924,9848,2227,4454,8908,475,950,1900,3800,7600,15200,12931,8517,
                   1737,3474,6948,13896,10451,5605,11210,5079,10158,2847,5694,11388,7355,14710,13999,
                   10525,5753,11506,7591,15182,13023,8701,1977,3954,7908,15816,16339,15333,13193,9041,
                   737,1474,2948,5896,11792,6243,12486,9679,4061,8122,16244,15019,12565,9833,2193,
                   4386,8772,203,406,812,1624,3248,6496,12992,8643,1989,3978,7956,15912,14355,
                   13413,11401,7505,15010,12551,9805,2265,4530,9060,651,1302,2604,5208,10416,5411,
                   10822,4303,8606,1919,3838,7676,15352,13235,8997,521,1042,2084,4168,8336,1379,
                   2758,5516,11032,4723,9446,3471,6942,13884,10299,5173,10346,5271,10542,5663,11326,
                   7231,14462,13503,11581,7737,15474,15527,15629,15961,14577,13729,12033,6721,13442,11591,
                   7885,15770,16247,15021,12569,9841,2209,4418,8836,331,662,1324,2648,5296,10592,
                   5763,11526,7759,15518,15743,16061,14649,13873,10273,5121,10242,5191,10382,5471,10942,
                   4415,8830,191,382,764,1528,3056,6112,12224,7107,14214,11087,4829,9658,3895,
                   7790,15580,15867,16309,15145,12817,8289,1153,2306,4612,9224,3155,6310,12620,9947,
                   2549,5098,10196,3051,6102,12204,6939,13878,10287,5149,10298,5175,10350,5279,10558,
                   5695,11390,7359,14718,14015,10557,5689,11378,7335,14670,14047,10749,6073,12146,6823,
                   13646,11999,6653,13306,9143,813,1626,3252,6504,13008,8675,1925,3850,7700,15400,
                   15379,15461,15497,15697,16097,14721,14145,10945,4545,9090,839,1678,3356,6712,13424,
                   11427,7429,14858,12375,9453,3481,6962,13924,10379,5461,10922,4375,8750,31,62,
                   124,248,496,992,1984,3968,7936,15872,14403,13509,11721,8145,16290,15111,12877,
                   8409,1521,3042,6084,12168,6995,13990,10511,5725,11450,7479,14958,12447,9597,3769,
                   7538,15076,12683,10069,2793,5586,11172,4875,9750,2159,4318,8636,1851,3702,7404,
                   14808,14323,11173,4873,9746,2151,4302,8604,1915,3830,7660,15320,13299,9125,777,
                   1554,3108,6216,12432,9571,3717,7434,14868,12395,9365,3433,6866,13732,12043,6741,
                   13482,11543,7789,15578,15863,16301,15129,12913,8353,1281,2562,5124,10248,5203,10406,
                   5391,10782,4223,8446,1471,2942,5884,11768,8115,16230,14991,12637,9977,2481,4962,
                   9924,2507,5014,10028,2587,5174,10348,5275,10550,5679,11358,7423,14846,14271,11069,
                   4665,9330,3239,6478,12956,8571,1717,3434,6868,13736,12051,6757,13514,11735,8173,
                   16346,15351,13229,8985,625,1250,2500,5000,10000,2659,5318,10636,5979,11958,6447,
                   12894,8447,1469,2938,5876,11752,8083,16166,14863,12381,9465,3505,7010,14020,10699,
                   6101,12202,6935,13870,10271,5245,10490,5559,11118,4767,9534,3647,7294,14588,13755,
                   12085,6697,13394,11495,7565,15130,12919,8365,1305,2610,5220,10440,5587,11174,4879,
                   9758,2175,4350,8700,1979,3958,7916,15832,16371,15269,13065,8785,225,450,900,
                   1800,3600,7200,14400,13507,11717,8137,16274,15207,12941,8537,1777,3554,7108,14216,
                   11091,4837,9674,4055,8110,16220,15099,12725,10025,2577,5154,10308,5323,10646,5999,
                   11998,6655,13310,9151,829,1658,3316,6632,13264,9187,901,1802,3604,7208,14416,
                   13539,11653,8009,16018,14695,13965,10585,5873,11746,8071,16142,14943,12541,9657,3889,
                   7778,15556,15819,16341,15337,13201,9057,641,1282,2564,5128,10256,5219,10438,5583,
                   11166,4991,9982,2495,4990,9980,2491,4982,9964,2459,4918,9836,2203,4406,8812,
                   155,310,620,1240,2480,4960,9920,2499,4998,9996,2651,5302,10604,5787,11574,
                   7727,15454,15615,15805,16185,14897,12321,9217,3137,6274,12548,9803,2261,4522,9044,
                   747,1494,2988,5976,11952,6435,12870,8399,1501,3002,6004,12008,6547,13094,8719,
                   93,186,372,744,1488,2976,5952,11904,6467,12934,8527,1757,3514,7028,14056,
                   10643,5989,11978,6615,13230,8991,637,1274,2548,5096,10192,3043,6086,12172,7003,
                   14006,10543,5661,11322,7223,14446,13471,11645,7865,15730,16039,14605,13913,10481,5537,
                   11074,4807,9614,3935,7870,15740,16059,14645,13865,10257,5217,10434,5575,11150,4959,
                   9918,2367,4734,9468,3515,7030,14060,10651,6005,12010,6551,13102,8735,125,250,
                   500,1000,2000,4000,8000,16000,14659,14021,10697,6097,12194,6919,13838,10335,5373,
                   10746,6071,12142,6815,13630,11839,6205,12410,9399,3373,6746,13492,11563,7701,15402,
                   15383,15469,15513,15729,16033,14593,13889,10433,5569,11138,4935,9870,2399,4798,9596,
                   3771,7542,15084,12699,10101,2729,5458,10916,4363,8726,111,222,444,888,1776,
                   3552,7104,14208,11075,4805,9610,3927,7854,15708,16123,14773,14121,10769,4193,8386,
                   1479,2958,5916,11832,6195,12390,9359,3421,6842,13684,11947,6421,12842,8215,1133,
                   2266,4532,9064,659,1318,2636,5272,10544,5667,11334,7375,14750,14207,10941,4409,
                   8818,167,334,668,1336,2672,5344,10688,6083,12166,6991,13982,10623,5821,11642,
                   7863,15726,16031,14717,14009,10545,5665,11330,7367,14734,14175,11005,4537,9074,679,
                   1358,2716,5432,10864,4259,8518,1743,3486,6972,13944,10419,5413,10826,4311,8622,
                   1823,3646,7292,14584,13747,12069,6665,13330,11367,7309,14618,13943,10413,5401,10802,
                   4135,8270,1247,2494,4988,9976,2483,4966,9932,2523,5046,10092,2715,5430,10860,
                   4251,8502,1583,3166,6332,12664,9907,2341,4682,9364,3435,6870,13740,12059,6773,
                   13546,11671,8045,16090,14839,14253,11033,4721,9442,3463,6926,13852,10363,5301,10602,
                   5783,11566,7711,15422,15423,15421,15417,15409,15393,15361,15425,15553,15809,16321,15297,
                   13249,9153,961,1922,3844,7688,15376,15459,15493,15689,16081,14817,14209,11073,4801,
                   9602,3911,7822,15644,15995,14517,13609,11793,6241,12482,9671,4045,8090,16180,14891,
                   12309,9321,3217,6434,12868,8395,1493,2986,5972,11944,6419,12838,8207,1117,2234,
                   4468,8936,403,806,1612,3224,6448,12896,8323,1349,2698,5396,10792,4115,8230,
                   1039,2078,4156,8312,1203,2406,4812,9624,3955,7910,15820,16347,15349,13225,8977,
                   609,1218,2436,4872,9744,2147,4294,8588,1883,3766,7532,15064,12787,10149,2825,
                   5650,11300,7179,14358,13423,11421,7545,15090,12711,9997,2649,5298,10596,5771,11542,
                   7791,15582,15871,16317,15161,12849,8225,1025,2050,4100,8200,1107,2214,4428,8856,
                   371,742,1484,2968,5936,11872,6275,12550,9807,2269,4538,9076,683,1366,2732,
                   5464,10928,4387,8774,207,414,828,1656,3312,6624,13248,9155,965,1930,3860,
                   7720,15440,15587,15749,16201,15057,12769,10113,2881,5762,11524,7755,15510,15727,16029,
                   14713,14001,10529,5633,11266,7239,14478,13663,12029,6585,13170,8871,269,538,1076,
                   2152,4304,8608,1795,3590,7180,14360,13427,11429,7433,14866,12391,9357,3417,6834,
                   13668,11915,6485,12970,8471,1645,3290,6580,13160,8851,357,714,1428,2856,5712,
                   11424,7427,14854,12367,9437,3577,7154,14308,11147,4949,9898,2327,4654,9308,3323,
                   6646,13292,9115,885,1770,3540,7080,14160,10979,4485,8970,599,1198,2396,4792,
                   9584,3747,7494,14988,12635,9973,2473,4946,9892,2315,4630,9260,3099,6198,12396,
                   9371,3445,6890,13780,12267,7061,14122,10775,4205,8410,1527,3054,6108,12216,6963,
                   13926,10383,5469,10938,4407,8814,159,318,636,1272,2544,5088,10176,3011,6022,
                   12044,6747,13494,11567,7709,15418,15415,15405,15385,15473,15521,15617,15937,14529,13761,
                   12225,7105,14210,11079,4813,9626,3959,7918,15836,16379,15285,13097,8721,97,194,
                   388,776,1552,3104,6208,12416,9539,3781,7562,15124,12907,8341,1385,2770,5540,
                   11080,4819,9638,3855,7710,15420,15419,15413,15401,15377,15457,15489,15681,16065,14785,
                   14273,11201,5057,10114,2887,5774,11548,7803,15606,15791,16157,14969,12465,9505,3585,
                   7170,14340,13387,11477,7657,15314,13287,9101,857,1714,3428,6856,13712,12131,6789,
                   13578,11863,6381,12762,10231,2989,5978,11956,6443,12886,8431,1437,2874,5748,11496,
                   7571,15142,12815,8285,1273,2546,5092,10184,3027,6054,12108,6875,13750,12079,6685,
                   13370,11319,7213,14426,13559,11693,7961,15922,14375,13325,11353,7409,14818,14215,11085,
                   4825,9650,3879,7758,15516,15739,16053,14633,13841,10337,5249,10498,5703,11406,7519,
                   15038,12607,9789,2105,4210,8420,1419,2838,5676,11352,7411,14822,14223,11101,4857,
                   9714,4007,8014,16028,14715,14005,10537,5649,11298,7175,14350,13407,11517,7609,15218,
                   12967,8461,1625,3250,6500,13000,8659,2021,4042,8084,16168,14867,12389,9353,3409,
                   6818,13636,11979,6613,13226,8983,621,1242,2484,4968,9936,2531,5062,10124,2907,
                   5814,11628,7835,15670,15919,14365,13433,11441,7457,14914,12487,9677,4057,8114,16228,
                   14987,12629,9961,2449,4898,9796,2251,4502,9004,539,1078,2156,4312,8624,1827,
                   3654,7308,14616,13939,10405,5385,10770,4199,8398,1503,3006,6012,12024,6579,13158,
                   8847,349,698,1396,2792,5584,11168,4867,9734,2127,4254,8508,1595,3190,6380,
                   12760,10227,2981,5962,11924,6507,13014,8687,1949,3898,7796,15592,15763,16229,14985,
                   12625,9953,2433,4866,9732,2123,4246,8492,1563,3126,6252,12504,9715,4005,8010,
                   16020,14699,13973,10601,5777,11554,7687,15374,15455,15613,15801,16177,14881,12289,9281,
                   3265,6530,13060,8779,213,426,852,1704,3408,6816,13632,11971,6597,13194,9047,
                   749,1498,2996,5992,11984,6627,13254,9167,989,1978,3956,7912,15824,16355,15237,
                   13129,8913,481,962,1924,3848,7696,15392,15363,15429,15561,15825,16353,15233,13121,
                   8897,449,898,1796,3592,7184,14368,13315,11333,7369,14738,14183,10893,4441,8882,
                   295,590,1180,2360,4720,9440,3459,6918,13836,10331,5365,10730,6039,12078,6687,
                   13374,11327,7229,14458,13495,11565,7705,15410,15399,15373,15449,15601,15777,16129,14913,
                   12481,9665,4033,8066,16132,14923,12501,9705,3985,7970,15940,14539,13781,12265,7057,
                   14114,10759,4173,8346,1399,2798,5596,11192,4915,9830,2191,4382,8764,59,118,
                   236,472,944,1888,3776,7552,15104,12867,8389,1481,2962,5924,11848,6355,12710,
                   9999,2653,5306,10612,5803,11606,7919,15838,16383,15293,13113,8753,33,66,132,
                   264,528,1056,2112,4224,8448,1603,3206,6412,12824,8307,1189,2378,4756,9512,
                   3603,7206,14412,13531,11765,8105,16210,15079,12685,10073,2801,5602,11204,5067,10134,
                   2927,5854,11708,7995,15990,14511,13597,11897,6321,12642,9863,2381,4762,9524,3627,
                   7254,14508,13595,11893,6313,12626,9959,2445,4890,9780,2091,4182,8364,1307,2614,
                   5228,10456,5619,11238,5007,10014,2687,5374,10748,6075,12150,6831,13662,12031,6589,
                   13178,8887,301,602,1204,2408,4816,9632,3843,7686,15372,15451,15605,15785,16145,
                   14945,12417,9537,3777,7554,15108,12875,8405,1513,3026,6052,12104,6867,13734,12047,
                   6749,13498,11575,7725,15450,15607,15789,16153,14961,12449,9473,3649,7298,14596,13899,
                   10453,5609,11218,5095,10190,3039,6078,12156,6843,13686,11951,6429,12858,8247,1069,
                   2138,4276,8552,1683,3366,6732,13464,11635,7845,15690,16087,14829,14233,11121,4769,
                   9538,3783,7566,15132,12923,8373,1321,2642,5284,10568,5843,11686,7951,15902,14463,
                   13501,11577,7729,15458,15495,15693,16089,14833,14241,11009,4673,9346,3399,6798,13596,
                   11899,6325,12650,9879,2413,4826,9652,3883,7766,15532,15643,15989,14505,13585,11873,
                   6273,12546,9799,2253,4506,9012,555,1110,2220,4440,8880,291,582,1164,2328,
                   4656,9312,3203,6406,12812,8283,1269,2538,5076,10152,2835,5670,11340,7387,14774,
                   14127,10781,4217,8434,1447,2894,5788,11576,7731,15462,15503,15709,16121,14769,14113,
                   10753,4161,8322,1351,2702,5404,10808,4147,8294,1167,2334,4668,9336,3251,6502,
                   13004,8667,2037,4074,8148,16296,15123,12901,8329,1361,2722,5444,10888,4435,8870,
                   271,542,1084,2168,4336,8672,1923,3846,7692,15384,15475,15525,15625,15953,14561,
                   13697,12097,6849,13698,12103,6861,13722,12151,6829,13658,12023,6573,13146,8951,429,
                   858,1716,3432,6864,13728,12035,6725,13450,11607,7917,15834,16375,15277,13081,8817,
                   161,322,644,1288,2576,5152,10304,5315,10630,5967,11934,6527,13054,8639,1853,
                   3706,7412,14824,14227,11109,4745,9490,3687,7374,14748,14203,10933,4393,8786,231,
                   462,924,1848,3696,7392,14784,14275,11205,5065,10130,2919,5838,11676,8059,16118,
                   14767,14109,10873,4273,8546,1671,3342,6684,13368,11315,7205,14410,13527,11757,8089,
                   16178,14887,12301,9305,3313,6626,13252,9163,981,1962,3924,7848,15696,16099,14725,
                   14153,10961,4577,9154,967,1934,3868,7736,15472,15523,15621,15945,14545,13793,12161,
                   6977,13954,10567,5837,11674,8055,16110,14751,14205,10937,4401,8802,135,270,540,
                   1080,2160,4320,8640,1987,3974,7948,15896,14451,13477,11529,7761,15522,15623,15949,
                   14553,13809,12193,6913,13826,10311,5325,10650,6007,12014,6559,13118,8767,61,122,
                   244,488,976,1952,3904,7808,15616,15939,14533,13769,12241,7137,14274,11207,5069,
                   10138,2935,5870,11740,8187,16374,15279,13085,8825,177,354,708,1416,2832,5664,
                   11328,7363,14726,14159,10973,4601,9202,935,1870,3740,7480,14960,12451,9477,3657,
                   7314,14628,13835,10325,5353,10706,6119,12238,7135,14270,11071,4669,9338,3255,6510,
                   13020,8699,1973,3946,7892,15784,16147,14949,12425,9553,3809,7618,15236,13131,8917,
                   489,978,1956,3912,7824,15648,15875,14405,13513,11729,8161,16322,15303,13261,9177,
                   1009,2018,4036,8072,16144,14947,12421,9545,3793,7586,15172,13003,8661,2025,4050,
                   8100,16200,15059,12773,10121,2897,5794,11588,7883,15766,16239,15005,12665,9905,2337,
                   4674,9348,3403,6806,13612,11803,6261,12522,9623,3949,7898,15796,16171,14869,12393,
                   9361,3425,6850,13700,12107,6869,13738,12055,6765,13530,11767,8109,16218,15095,12717,
                   10009,2673,5346,10692,6091,12182,7023,14046,10751,6077,12154,6839,13678,11935,6525,
                   13050,8631,1837,3674,7348,14696,13971,10597,5769,11538,7783,15566,15839,16381,15289,
                   13105,8737,1);
constant inverses : numarray := (1,1,8737,15422,13105,10283,7711,13697,15289,4991,13876,12792,11566,3706,14561,6169,
                   16381,13366,11166,1182,6938,16129,6396,1494,5783,14076,1853,3797,15953,4264,11821,
                   3241,15839,1127,6683,6355,5583,10392,591,3992,3469,658,15777,4692,3198,1459,
                   747,1804,10602,4581,7038,12243,8639,906,9547,10003,15625,16243,2132,6214,13623,
                   7074,9333,10558,15566,6378,8210,14983,12076,11148,11848,13663,10438,16055,5196,10512,
                   8966,13315,1996,2596,9447,5067,329,13154,15601,6833,2346,3006,1599,8496,8440,
                   1443,9044,739,902,15687,5301,6621,10963,989,3519,13424,13768,8924,13054,14665,
                   453,15489,12420,8561,12712,9289,15525,16069,15768,6525,1066,891,3107,16208,14522,
                   11973,3537,398,12315,12813,5279,2751,7783,14932,3189,1651,4105,5744,16226,4603,
                   6038,4274,5574,6723,5924,15547,14478,1329,5219,11339,15738,10626,2598,13546,5256,
                   1687,4483,5424,14368,14537,998,1205,1298,297,12370,10989,11204,13450,8837,331,
                   6577,5743,15449,8821,12153,7724,1173,12629,1503,5072,8510,8198,4248,8187,4220,
                   8574,8432,7983,4522,5647,9040,11014,451,5247,15490,13760,10363,8558,11983,13415,
                   14152,5757,9167,246,9470,4917,6712,5732,6884,11843,4462,9541,6527,1564,16005,
                   4654,8899,9322,15457,12224,6210,12320,12953,10668,6356,6384,12293,6699,15475,10492,
                   15683,6847,7884,8014,11935,417,533,1437,9116,7952,9264,865,8104,5442,7261,
                   4062,13635,3769,9417,11551,199,9166,14892,15019,15143,3816,10350,7431,10110,13742,
                   11538,12123,7466,3531,9243,1243,8472,14140,10789,10105,2872,10840,8113,14745,10972,
                   15250,3019,15361,2137,1354,2787,1431,12032,10552,2962,7866,15484,7578,7239,6317,
                   8377,10036,10256,7892,13316,6228,7869,2453,5313,7986,1299,159,6773,13887,2628,
                   3996,8554,14075,10976,12543,2712,12721,7184,3396,15941,15646,499,16245,8315,16202,
                   649,2800,8885,10300,6185,15151,14167,8987,5602,5085,6725,6595,13155,82,8836,
                   165,12025,4356,10518,12778,15373,7363,13083,2448,13725,1790,3862,9728,8299,10888,
                   14987,13010,8398,3548,2536,10480,4255,13784,4099,5587,2124,13139,11740,2128,2110,
                   13009,4287,11297,4216,9381,11702,5466,2261,745,10534,15925,4520,3610,5507,16285,
                   8896,9857,10270,9780,7745,905,6880,7206,13852,6944,4279,10765,13638,15888,14354,
                   836,7076,13160,10527,10865,13254,12578,123,3536,4735,16174,11195,12218,3356,9263,
                   2866,5225,3442,6774,13568,13231,2231,2497,12419,2265,11934,231,782,16265,15715,
                   11429,2327,915,13120,2370,4661,12497,15377,11142,6112,5564,3105,6073,6160,10232,
                   15213,9407,5334,10498,3178,15948,3192,1957,14883,2134,12084,5030,15384,4928,5246,
                   188,15488,106,12158,12308,3942,4652,4007,12740,13678,6402,8945,15184,9003,13002,
                   8431,9155,4558,2729,3976,13210,4632,2789,9105,5273,4052,2008,2721,7978,11279,
                   16351,2031,9626,14464,4998,9597,12546,12357,12772,13486,7250,8770,11515,4583,15608,
                   7446,3760,16244,312,16306,3939,1908,11506,5175,14533,11426,8722,5055,13861,6871,
                   2385,5769,15118,13708,5900,3733,12316,9412,11810,12332,7345,8268,11138,4236,7694,
                   7070,2912,14131,15743,12701,1424,1436,232,5420,15172,11769,7086,16109,13723,5486,
                   10786,7625,1313,10180,16355,15393,10612,9741,8375,677,15277,10064,4350,8426,14740,
                   6016,15285,5276,3714,1481,10345,3933,16383,7742,2976,3789,7081,11266,7375,11895,
                   11421,12925,3022,5018,3931,5128,15308,3946,3776,6658,15445,3114,5903,11647,4108,
                   9963,13949,10305,6657,3993,38,8360,10993,8814,2411,12059,6887,14654,2302,1314,
                   16032,1998,12837,4277,4284,14684,14299,5488,2790,14942,4013,1356,16051,15097,16009,
                   3592,7448,1698,14946,15619,3191,7823,15886,8920,7521,15771,11655,12828,8832,8101,
                   7083,9061,4470,1400,14423,13179,15985,5150,1639,11829,4608,16310,13601,14730,6651,
                   13228,12742,2801,316,11215,10906,12035,7643,11968,5616,15248,1200,41,3468,4418,
                   2924,8819,11487,13661,7252,2178,11545,5259,9710,6389,11944,15399,1975,11328,3635,
                   15276,550,1224,15230,14575,12499,895,2514,1931,4453,4864,10376,12820,11288,5444,
                   5402,16228,6806,6505,4223,4199,3111,1774,7791,1268,11814,5240,8228,10862,12963,
                   6892,5541,10784,6127,10440,15347,1062,6174,15240,5572,5870,16034,1064,16300,1055,
                   1457,15177,12630,10878,8553,13361,11525,2108,6398,12403,2644,5851,10881,2733,8276,
                   9803,14242,9045,93,5267,10566,15675,4758,2260,369,1805,46,10464,10051,15855,
                   10146,4448,3220,12641,7852,5135,3734,4890,9539,11521,5396,9189,1854,3440,4175,
                   3603,3117,6926,6814,3472,6857,10874,1209,14119,11210,6819,11989,7944,14408,7177,
                   12876,418,16264,3538,5774,6580,13349,13998,4025,14105,6007,6627,11218,6289,8470,
                   8732,6600,1768,1569,11038,8493,8087,5650,14332,3012,6109,13402,1678,5364,12342,
                   13911,1433,2934,10261,7540,1721,1529,3387,10302,6784,16135,15350,10188,9850,6376,
                   9921,1941,14944,16154,9805,16204,5967,6164,8786,16029,391,14355,15845,1616,15504,
                   10043,13427,10514,9898,10503,9192,7515,6560,1236,1185,4181,11067,11438,14921,1363,
                   15401,10443,5571,5422,3056,3214,2782,14589,9265,237,10749,2636,3080,13325,5116,
                   5346,16279,2798,12414,3482,2667,11217,5249,1907,1589,11880,7974,1918,1596,12835,
                   8691,1396,16176,11689,1067,117,6042,4629,2515,682,7692,3042,2464,11889,2623,
                   13739,94,15686,7744,381,53,8638,6079,7660,6154,3098,1971,3757,2326,423,
                   9714,10706,6370,1295,6839,10570,3201,10471,13145,14867,7592,1526,13236,14648,6501,
                   4936,12886,3249,13248,4090,2279,15345,10101,7880,1988,13393,6605,4401,2316,12535,
                   10067,10979,13289,7408,10349,7267,2026,10496,1004,11662,10097,10206,3989,1766,13350,
                   4846,15822,5861,8662,8904,4813,4215,7232,13440,2499,16263,12447,15439,6273,12938,
                   14851,4262,6386,6986,6743,3570,3625,13117,4385,7512,13404,15375,10962,99,7804,
                   8794,3723,6224,1880,14123,8122,7068,156,1204,8153,3739,9616,9657,954,11663,
                   5753,9685,10298,6309,15939,14208,5713,1904,4361,3957,11262,8641,14643,12435,12106,
                   10489,9865,15979,10597,5593,7559,2340,6854,3766,2950,6231,9579,10269,6158,9086,
                   4706,4209,5905,7667,6166,13680,11385,2147,4134,4736,5569,10404,2118,14610,3847,
                   1793,3535,1995,1456,720,14776,7162,15518,2096,15087,11992,712,6175,718,16301,
                   116,890,2710,1719,7586,2420,13533,7347,3543,14064,15703,16194,14572,10052,2743,
                   6859,5393,1417,11461,7319,8369,14592,5090,1332,15824,3674,15409,3491,5306,5101,
                   12583,13292,12922,10069,9075,12990,16375,8825,5032,4486,2175,7297,4213,4323,7370,
                   10244,3008,7720,16379,4992,2638,5501,1857,6619,8389,7734,13845,13997,9615,7491,
                   15838,33,3871,9844,1488,14089,9543,5125,12277,1263,5633,5212,11334,13219,13594,
                   13575,13423,10622,15135,11562,1511,3927,2509,6768,9612,1198,2564,12694,7654,15007,
                   1973,6703,1888,8141,3329,5314,15371,1828,1557,3973,10662,12120,13470,14391,2054,
                   16122,12628,172,14623,14181,13825,15807,12065,15594,9709,8042,19,11167,4180,850,
                   14169,16012,4407,12256,9876,10800,13740,10033,12114,6342,7327,6237,1151,9613,657,
                   15249,8016,1435,999,157,15155,15748,10875,773,2142,7170,7342,10755,14796,9359,
                   2744,15971,1395,9267,7471,2566,9719,7498,678,15231,15736,9409,16221,7034,15717,
                   10813,1796,11929,3724,11372,849,6561,7473,1657,15520,14304,9242,261,11622,11268,
                   7943,14225,4460,15183,11409,11049,15596,13049,13538,12479,6414,1366,4416,9038,11763,
                   8158,12276,1135,13203,13102,2235,10398,700,11815,15882,5071,15260,14948,15641,5807,
                   2575,13945,8466,3480,13627,7582,2304,2442,8155,13702,14513,10419,7365,6470,11996,
                   6101,6614,11840,6371,919,10073,5496,158,296,14278,9973,5453,4548,13728,5680,
                   11468,9842,5984,11257,2808,12055,7624,543,600,16033,8757,9385,1734,2232,2209,
                   2517,1462,6478,13080,9011,13390,4870,14479,143,3626,12731,1089,5091,13485,9433,
                   10340,3373,4855,16087,11867,3236,5972,14678,15410,10501,8698,2313,5664,3044,9528,
                   10551,7638,13758,275,2136,612,16050,7615,11327,15958,2760,14920,855,9118,9259,
                   1257,6415,8676,7492,10899,13716,2432,14045,5188,10556,6410,14228,5644,7963,2722,
                   12751,2701,4765,8114,12279,3403,7340,11925,15658,10782,1724,10770,2860,9266,1218,
                   887,8690,11542,1746,634,14422,5907,12397,2620,11788,4114,13198,5431,15783,15216,
                   5512,3446,16338,10483,12850,5392,1083,10710,7015,5220,15378,16344,1875,531,12700,
                   3087,9753,7620,16107,2786,277,2935,812,8017,1203,532,233,8150,4577,8238,
                   3991,8441,91,16261,14853,6315,2345,5439,3166,12949,10678,14393,6241,13475,5115,
                   1054,721,3199,45,14872,9281,1322,6479,10572,15353,14177,1626,10103,14519,4138,
                   4541,12548,4639,7121,2060,13195,5515,8719,16076,10344,560,5283,11578,15548,7048,
                   2379,6129,1130,14088,8857,14376,8615,5368,23,6397,5232,6821,12672,8488,15574,
                   9423,5073,174,2224,6059,1610,14213,14993,15427,3926,1146,10278,12648,1867,9336,
                   2445,12507,12416,15789,13473,1794,2698,16269,13267,13298,927,7593,1720,817,10758,
                   13969,9512,11356,9271,7066,3463,14178,3407,5882,1736,3332,12101,2163,5437,6686,
                   8317,14341,14770,1822,5605,11317,12144,15073,13643,8396,3972,1164,7204,13883,11301,
                   9137,6438,14254,209,6526,8132,9436,1769,799,2887,8717,3290,11620,14387,9695,
                   6999,10346,9725,13659,14765,12104,10650,2898,11984,15136,5609,5333,11881,880,4235,
                   13669,4366,11005,3300,15943,884,12834,8497,88,5519,14600,12983,8634,11754,5106,
                   2825,1722,7166,13185,1506,14212,10703,7051,6701,7637,839,15844,2682,6183,6171,
                   5461,14602,13689,8429,2407,1467,14176,13867,16275,3770,15009,8573,5649,8413,10592,
                   9404,9453,5151,639,3392,5787,15778,3417,7675,3144,5094,9132,4925,14783,3188,
                   131,12609,10690,8683,5779,7472,1239,8077,4010,12551,11085,8102,11727,10630,15900,
                   3082,2081,4393,11966,15727,10734,8930,14434,15912,13075,15571,6093,808,5365,7752,
                   9035,12732,14110,14360,7037,5257,151,4949,13656,13986,2691,4596,5181,11404,8769,
                   3280,8727,618,14947,8305,14682,10763,11766,14268,5511,5719,13512,16133,12291,8328,
                   5521,15413,5626,13892,13222,10432,2093,2711,1069,1528,816,1607,2824,1391,10783,
                   15967,8827,12345,2439,8791,10885,14047,14721,1318,2233,1540,3333,14375,7203,2558,
                   1750,2673,5171,15850,15395,1399,11543,6207,12407,1741,2559,10004,14699,14281,13253,
                   10337,4651,8600,11425,8507,11912,5940,13110,3987,14934,959,3988,798,1568,15152,
                   10657,13016,4579,698,7790,8088,6906,13557,6575,8244,15128,8731,15074,3021,1962,
                   11051,13429,9928,8633,341,13724,3846,1051,1521,13472,1232,11928,13593,4037,10046,
                   6232,14580,12493,47,746,7843,10333,3872,9933,8863,14413,8763,2660,4319,16252,
                   10750,7361,3830,13343,3077,9351,1549,14771,8696,12808,9591,4766,1163,15370,8946,
                   7432,4857,3698,5353,5548,3185,2182,8358,6338,12154,8543,5285,12613,9313,6491,
                   13906,8448,15245,3666,16168,15598,3796,26,763,9188,6618,1118,7324,11680,11923,
                   12450,2468,4761,6443,10896,9337,1514,6624,16304,2045,12644,9810,5476,16345,1423,
                   12699,2937,3940,5534,994,14122,14345,2058,11975,3260,10937,10633,1158,8140,14938,
                   14248,12680,8703,14160,9662,15317,4914,3704,13419,13847,14861,11280,11629,1013,5712,
                   5248,879,502,11507,5831,4982,12697,6915,5103,3636,9707,2883,883,7975,6675,
                   13163,2423,3584,7911,4895,10579,15070,4331,11395,4452,684,11079,4422,10778,2217,
                   3616,12433,6720,14012,9920,827,15842,2889,14958,9340,15366,15573,11873,9655,6469,
                   3960,16160,9817,2131,15862,3193,443,3493,8347,12042,13977,1785,3020,9525,10038,
                   15295,9808,10929,15141,3756,912,6702,1156,15398,673,5481,7093,8720,13243,3902,
                   8595,4397,15077,9572,9181,3112,14302,940,13392,14772,9763,4061,12525,3534,1053,
                   78,2597,602,12836,11725,2569,9580,10185,4808,3318,12541,16288,477,4053,13542,
                   10857,10525,6758,12491,13747,5149,6973,11891,16044,15616,14800,7104,7729,10505,10987,
                   952,10497,10917,13125,9627,482,5631,6264,12993,7556,16056,12604,14952,3875,6053,
                   3163,13917,11376,12645,1870,15636,14511,13971,11172,10445,5254,11490,8642,1170,16123,
                   3427,2812,1883,14344,1475,7120,11786,11336,12436,14084,13871,2088,3079,2940,4543,
                   15870,2353,14624,10777,15001,10665,2805,11480,11477,3083,1667,6840,13610,13341,10661,
                   9744,6882,2067,13870,2368,8860,10433,1717,5202,11121,1059,15519,7305,6220,9634,
                   13004,8609,11522,9414,6141,8644,9624,728,6399,360,13008,7388,9642,3581,8842,
                   7759,11915,1048,14611,16214,7649,5996,9466,356,13138,11822,12273,359,11741,15863,
                   1954,58,6215,445,14882,1355,274,8570,4187,3793,16330,1210,7171,14415,12112,
                   11384,1043,9418,15058,7032,13795,15498,8162,8097,14706,7286,9702,5026,15033,10106,
                   8424,12100,1543,10409,7495,8421,14031,13379,5472,11370,15201,12921,6691,7296,1106,
                   2545,7631,666,11544,7912,14785,1837,3184,15417,5706,9456,13035,2653,6694,11223,
                   3829,15026,15270,6646,6191,6461,13381,12683,13059,13208,7901,6495,7041,15834,15781,
                   13085,3455,2516,1320,2243,3866,9758,13383,11361,8364,10779,1935,10832,8213,3685,
                   10354,5122,10137,1504,6058,3860,11342,15836,11861,2496,412,1319,1735,10399,1266,
                   8577,7938,11980,15656,12867,10850,3867,2210,14635,3801,14711,8049,12518,2399,11392,
                   13650,7919,4457,8753,12711,9646,9894,4922,5859,744,368,14757,14832,12418,415,
                   10275,15751,13787,2771,8278,16317,10529,7647,2606,8694,5667,10387,15344,936,6797,
                   8073,14498,6588,14358,11058,5311,15528,16302,8689,5781,15793,8402,15556,9610,7442,
                   9927,7420,3384,4727,4806,14981,599,14655,1282,2443,6347,16328,3827,12193,16238,
                   8095,8699,1347,12086,3229,944,12534,11719,9801,9377,9226,2657,15975,15396,5251,
                   914,422,8491,10292,9699,13321,5331,11386,6060,7780,6735,11088,15930,15918,1027,
                   7558,8061,7293,6314,1447,86,3007,16046,5109,14739,6544,14625,2072,15614,7611,
                   13745,11258,7797,6268,12503,10517,4021,6770,8744,11310,14318,14877,2090,8861,425,
                   13121,14733,13466,8006,15415,10938,13497,6128,1486,4938,5210,5400,3654,6870,511,
                   12729,7989,6057,4291,3171,7569,11374,7936,11791,8008,8222,13537,12519,2249,9065,
                   6937,16361,4600,4008,12875,8428,1625,9170,14137,8815,595,16312,5890,7874,5126,
                   14108,13439,9123,5078,1071,7587,3585,1922,3671,2775,14112,14831,7398,12453,12390,
                   6573,1372,14044,15632,2654,8344,5721,12344,1729,11446,7561,1283,2305,12506,1516,
                   3749,15820,339,13082,16286,12785,7868,293,12353,6974,15759,3794,3517,4301,15507,
                   4516,14143,10128,898,11888,13677,13957,1862,4760,5686,4785,9097,8363,12017,14786,
                   11449,6587,8477,8021,7760,10010,7152,15492,4621,8118,8867,10810,5811,3147,5634,
                   3822,11682,5081,14825,13107,2230,413,16262,970,13417,7008,14261,3573,7798,3703,
                   15197,14290,6769,1148,14974,11359,3207,4316,683,894,2208,1321,4519,10577,13528,
                   8617,4079,9649,6138,16231,8214,10251,15336,6279,6551,7129,9852,3471,5199,14421,
                   350,10481,13618,4838,7941,15303,11206,11457,7630,2176,7474,3292,15533,16196,10614,
                   7274,10022,3210,14621,13942,4233,11527,1740,1751,14524,4444,3791,4830,1152,12695,
                   1221,7470,11724,2001,6851,11111,15993,9316,13944,1276,11331,10194,3235,7923,5998,
                   7395,10699,16075,3307,5344,5920,13771,11856,11202,9194,6118,12685,8309,2748,14583,
                   79,1997,148,13547,7139,4188,12635,8878,10375,4762,2274,8695,6864,7383,2840,
                   5727,5734,9093,4921,15465,2992,11816,14301,12066,1404,11789,13738,900,3812,15369,
                   9006,4102,300,3997,15729,11743,13115,5837,12405,6571,867,10748,1116,5500,9841,
                   7733,9931,5856,731,12402,3239,11827,6540,4899,13240,13128,6695,2188,2435,15633,
                   15974,2322,8806,15668,1813,8762,15100,4773,8193,7349,11216,876,14455,14503,12365,
                   10013,5170,1742,9399,8046,11098,11529,15690,9977,13580,10006,1618,6182,2986,12040,
                   7339,10548,7705,6981,13987,1691,4349,3649,9893,6459,2832,5478,1522,16268,4764,
                   1382,14010,14677,3819,13401,6879,11092,8872,15424,1068,1718,306,12720,8025,16143,
                   11518,12817,13374,6334,7979,478,1380,12750,7460,9441,9098,7454,4559,469,12340,
                   11589,8277,734,11942,7259,4338,8869,3746,5394,14184,12885,6858,1080,1216,15970,
                   14671,3465,2594,14582,5278,127,3205,15227,7114,11065,2822,9047,11692,13905,1361,
                   15959,15046,8250,10087,14056,11119,3758,4057,14194,13786,2269,9348,10828,3670,2425,
                   13675,10871,7829,4479,5391,11965,862,14588,5385,10846,1430,276,4633,473,609,
                   5489,9114,8196,4345,15132,5771,12001,873,16278,317,648,7211,10397,10664,2077,
                   14871,11640,1310,12054,5894,16019,2057,3426,6599,12530,10426,4980,15602,4411,7608,
                   7927,2756,9046,1723,1606,8169,16039,13912,5075,6425,12786,2696,5479,8252,13719,
                   5355,13476,12178,6132,2610,5726,7689,4940,8172,6067,8584,10953,9000,16060,6350,
                   6776,9254,4370,12589,12638,3810,14669,15700,11729,1393,10771,8875,5682,10138,13851,
                   406,5224,11657,15330,8312,13152,266,10841,8789,15905,4075,6303,10961,3547,4119,
                   7173,9706,1917,12893,6531,8716,1570,15843,1943,16163,10681,11892,6786,9909,6015,
                   10430,3089,1583,10651,15211,13131,5339,15987,15933,6292,11793,14530,14448,3041,11228,
                   6363,527,7071,9033,9966,9246,15980,8759,3609,7436,6997,12289,11032,661,4419,
                   11910,13093,5286,9846,16349,10272,14737,6925,813,1432,12698,1877,15994,7826,2069,
                   3078,11007,4141,6274,4826,11054,5620,12233,15326,1030,6230,15332,9371,10468,12960,
                   13094,3143,8038,6762,5172,3155,280,7867,10352,15281,5789,12666,7774,7810,3524,
                   6110,9860,11568,10713,11634,565,7743,7044,14760,13165,14441,7188,12330,13042,9506,
                   2684,12041,8746,14912,11871,4219,2616,11817,12147,8952,6336,11979,4244,5160,7787,
                   15436,12358,10867,11209,5659,87,2347,1112,7721,10740,4777,805,14333,14819,6645,
                   16233,8177,15360,272,1963,1784,573,12924,5139,8648,6324,12439,8580,4450,4668,
                   12301,9959,16346,14924,9146,6208,4529,15607,15322,14449,2909,897,7693,1349,5665,
                   15847,10025,15304,6994,6649,9673,9198,12388,11509,5942,860,3215,9145,5182,5379,
                   12162,14697,4097,4756,12904,5678,12476,12346,5048,3533,9215,9442,11499,7089,3255,
                   9350,1820,2941,2068,868,13324,1666,2080,13699,10920,9752,1426,10431,2897,3343,
                   5366,12831,8331,15907,13294,7385,12212,911,6155,10451,8939,13371,9391,6072,432,
                   16209,118,14468,8256,4198,697,1986,14303,582,5902,3602,767,14652,12268,13363,
                   14803,13305,12049,3219,15328,7127,6950,8777,9309,3263,16240,4066,10797,4718,12865,
                   8533,5888,9134,13201,10114,13063,13095,2957,1645,7674,5810,2489,15928,16198,12494,
                   8148,12170,5843,5173,2961,12511,4688,14476,9897,16119,7484,6052,2041,5325,7551,
                   1449,5438,5992,3678,7568,2390,10453,15313,10315,5700,13589,13364,440,15949,10852,
                   5113,14483,6728,2183,1836,14175,5885,1650,130,15618,621,442,1956,6417,10586,
                   12985,15639,44,1458,10470,922,7300,3245,15226,2752,4317,2512,5877,7996,2553,
                   10023,10149,14604,861,3057,3583,6863,15329,3124,753,4449,7106,8779,14022,9451,
                   12260,15672,12087,2315,11467,12092,9090,13412,7922,2578,1341,11866,11826,2646,11820,
                   31,10379,14014,7301,3203,14493,14080,12887,933,9874,8404,8444,13232,7088,3075,
                   14644,16150,15848,8685,1885,11974,16241,3130,12959,8443,10537,16173,12879,14839,5296,
                   13816,4702,12954,12375,14256,10286,4033,8990,14496,1696,8726,10604,15093,7889,9387,
                   9357,11691,11484,11171,1572,11621,2547,7475,4566,6277,11199,13448,16126,9637,1594,
                   15942,8800,12522,14977,14330,5345,2584,13012,3712,10600,12934,3736,5093,8266,13123,
                   11751,14270,2005,4809,15010,9277,14215,4388,4051,14165,13510,4001,5315,1160,7950,
                   12324,1541,1737,9777,11798,10933,8855,5983,10781,15510,12708,5367,3090,4465,8371,
                   7217,4378,7956,9291,15272,3944,15432,12932,10695,11230,404,9262,10331,6685,3876,
                   11150,13188,5829,6366,9510,7055,4833,7180,11348,12191,7142,10341,1337,8810,11670,
                   11147,16356,6828,4026,6993,5918,10080,13963,2298,4726,10303,818,5702,8955,13057,
                   7606,1640,5786,13098,10720,309,7185,16144,14964,12825,14087,7341,1386,14116,8623,
                   5883,1538,7134,6635,10466,13558,10506,12746,6756,13591,15779,1643,14880,5845,4164,
                   8318,10473,16071,15419,4751,2813,2056,6946,5484,6611,7164,5216,11594,9783,4768,
                   10090,15554,8247,4841,764,4174,408,6775,8450,10213,1412,16339,8342,15894,14126,
                   6679,15630,3554,13084,2207,14909,10099,9954,11443,13066,5749,14179,1536,14670,2747,
                   16097,7354,659,40,9853,2533,770,6856,9379,6254,15922,9325,11312,14658,1279,
                   8467,875,12415,10009,16093,10296,4910,7925,6517,15408,1093,8346,1958,13482,14055,
                   11838,6098,14874,5269,8519,10343,9950,7756,5002,5363,16020,6125,14789,10647,15299,
                   9732,13841,12002,11060,7899,4300,2458,13425,100,12988,8260,5956,15517,2970,6111,
                   6555,9664,9704,13616,7467,259,9214,3070,1994,1052,399,122,784,5775,7576,
                   16200,14065,1074,6508,10429,10960,2879,349,8399,3895,15434,4044,6444,3453,15631,
                   14427,5508,12022,4863,4122,9681,7564,13902,13100,14288,7537,6816,10183,8378,981,
                   6742,14260,2503,14363,13322,4964,11715,13053,8494,8843,2114,6862,3216,1923,2422,
                   8236,13926,8409,15192,6736,10229,616,7449,5964,15662,14509,11854,9667,9395,5023,
                   13327,3116,766,7290,5499,14919,16299,8758,2919,373,4521,11632,11962,13839,11631,
                   1936,12432,12615,12632,13166,4739,15879,4289,13116,982,1330,12730,10830,6413,8126,
                   10240,5375,5275,11329,675,1915,5102,14382,4169,9251,4137,12386,4312,8487,7208,
                   16120,11132,4348,2693,6404,12852,12442,15301,2383,5401,8292,10629,7685,7627,4473,
                   13024,3716,12472,11101,12654,1849,15244,10325,5673,2774,2424,9241,11771,1091,15825,
                   4179,6934,3169,5993,6077,15451,12942,7849,10355,2220,14979,7237,12305,11009,11916,
                   13730,6953,7960,4224,6889,16359,11998,1833,4856,8084,11225,7799,2505,1898,13418,
                   13,11567,9052,10793,4594,12393,3309,13013,559,5277,3662,12473,5840,4985,13672,
                   4590,6225,992,1234,11373,11117,5454,11956,16112,5448,12136,12317,516,757,5134,
                   3312,5092,8152,1001,8671,13596,6322,16003,4905,3935,2738,5395,15821,2446,8422,
                   15462,15084,3825,10141,15653,1970,913,2767,11118,497,7447,7061,11445,15909,7671,
                   1029,6855,13634,243,1630,15008,14205,11570,14053,10648,579,3947,4070,4682,7469,
                   9050,7124,11180,6340,8774,13022,10902,7080,566,4831,2562,16331,2140,2457,15758,
                   1852,27,14356,5001,14634,2245,16167,6782,5640,15805,13463,7231,9179,7915,2856,
                   14668,2624,15368,9110,5088,251,15142,13400,2704,10562,6727,2491,5635,15085,3753,
                   12192,2308,11222,2191,1818,13342,12500,11808,10112,14347,9112,6290,11698,15832,12072,
                   15859,15252,14155,9882,15175,1792,1050,11602,9296,11182,15710,13960,5039,7535,12099,
                   10836,15692,13408,12004,2226,11343,342,9729,14210,13277,2211,2242,5389,12658,9845,
                   1128,1808,9932,14953,2039,3360,11151,7006,6487,4960,14293,9148,12753,7921,8687,
                   10117,5936,7479,9172,4670,12521,7683,15577,15435,3550,13585,13181,12538,5008,11907,
                   14729,1980,8594,8080,5938,12557,16340,9736,8184,7931,14429,9245,5878,8956,14554,
                   9459,10636,12908,11441,6021,5371,14701,15428,8541,11432,1510,1147,12475,8310,5019,
                   575,16382,562,4904,3745,14201,4828,16307,501,1878,5535,456,4653,3351,15273,
                   578,3777,7699,4649,9073,7271,10389,12995,12283,9788,4360,1015,15356,8912,1951,
                   6468,13032,15218,10935,13563,16211,10369,4786,4474,13263,11107,1556,1165,7151,6660,
                   470,13211,6696,11251,7386,11290,12592,9751,9679,14521,14935,1764,1767,958,8239,
                   1441,39,590,10035,11668,301,2629,6418,9071,13511,3327,10021,4748,4790,14024,
                   12741,458,2404,12874,1659,8076,14943,611,8144,11396,8911,15957,9675,5916,6771,
                   2362,14101,5350,13999,789,3379,6829,14916,14245,14584,4713,10287,3277,12223,9410,
                   13592,1799,8022,4697,7808,6381,7400,11302,3552,6445,11577,15005,13989,10196,14164,
                   3324,476,2009,13985,10671,14195,2768,15235,4970,12524,1992,241,7260,10462,9429,
                   3132,10796,15169,7907,3778,4683,8028,9174,6302,2876,7476,12109,9648,2522,10739,
                   4306,9228,14969,14607,15628,5688,10242,14995,13508,935,13249,7818,8498,15990,7193,
                   14696,3063,5586,354,13895,10390,2627,9007,5745,132,4321,5052,585,11646,15708,
                   4792,9360,9503,1406,13199,8588,10774,7172,2880,8384,9279,3560,9680,5893,5526,
                   5668,10437,6218,12651,7042,8306,14646,6628,1044,4737,9250,3641,1470,4540,11006,
                   2943,7935,13920,9913,15223,7312,13798,14125,4433,16237,9978,14069,8262,10075,7858,
                   5740,15061,13387,6842,9252,11354,8544,14458,3420,8319,6805,11382,14383,3639,14067,
                   6896,4872,6984,3441,765,9768,10826,6935,3676,1184,851,4430,13530,13889,8928,
                   8571,2139,2601,7138,14233,10653,8240,14325,15470,7047,11365,10167,3110,696,4817,
                   4584,6502,14961,13041,13031,5761,10795,4707,1037,10719,7500,4322,1108,4812,967,
                   364,9380,11870,2991,180,8575,6504,695,3694,6888,4821,13079,9439,6433,4421,
                   9793,11526,2556,13668,1590,524,7695,16040,16314,8107,8652,11473,14418,2998,5161,
                   4733,7158,178,8186,6569,11592,5911,6481,13785,352,8850,8932,13519,5263,15578,
                   10236,977,14850,29,15952,11778,15867,8959,10061,7441,6837,8324,12094,137,6039,
                   4285,604,10764,386,9545,16222,8165,4615,605,4276,11296,362,15878,3623,6056,
                   2389,5692,4667,8232,11938,4709,7806,7529,15666,3516,2459,14544,14559,7749,16148,
                   4081,10738,11761,12597,7353,10761,3643,12387,4851,10059,2513,3206,16253,1814,5053,
                   4106,4212,1109,6050,12869,8482,6665,13941,15495,11394,1928,12883,15500,14662,11897,
                   14336,10173,2736,8868,5685,11556,16273,15840,15133,2794,12080,4550,3648,2692,553,
                   10065,9945,6585,11462,10384,333,12024,5772,14809,3956,1014,16065,6562,8631,12677,
                   1592,11004,15421,6849,2853,9255,4728,5976,15188,12964,9999,15968,3347,7216,14282,
                   5322,9563,11390,7513,984,7635,7570,3323,14214,11830,11503,11967,1668,14339,4427,
                   15076,1982,15264,6781,6604,943,11599,5316,11918,6748,12257,1188,7917,7679,15603,
                   2819,15279,14591,9374,7109,1258,9039,660,2925,9792,4230,1933,11078,4879,8512,
                   14338,4395,13329,12977,4182,13531,14124,4149,8678,8845,5416,11366,12843,5206,9491,
                   14475,5177,5929,2561,14525,12781,10358,752,3221,3029,8581,1930,685,5671,14571,
                   7918,2253,13579,16165,1248,15182,206,9540,8370,3344,8514,14144,13934,5607,633,
                   9060,13025,3660,3969,4787,5990,11406,7828,2779,15104,6271,5425,152,9644,9208,
                   1105,5033,16052,14049,9549,13565,16026,10991,11673,6556,6259,12302,9870,11648,5696,
                   8661,6825,5252,11606,8817,10901,14856,13113,10983,15090,15724,4823,8969,4947,12917,
                   2461,15506,10576,2518,372,3611,184,5646,16115,7562,7416,12468,6209,3037,8942,
                   4995,13872,15354,15586,12838,14540,8509,10056,10918,4139,1471,15871,2070,14001,6464,
                   11470,12591,1303,5452,4347,12081,10544,6091,13928,7628,7672,5584,468,2728,12135,
                   10158,11749,13029,7249,6559,3294,6276,7179,7597,5529,12691,10366,6070,7764,12789,
                   8151,1439,13017,1773,10603,49,15609,494,4201,4816,7778,8146,4805,15828,3721,
                   13673,12610,14813,3710,12392,1692,5180,11034,6104,2403,16360,16227,135,8970,13775,
                   16062,7064,641,11828,9956,15123,11844,4642,8164,4283,9560,7507,13809,11619,8119,
                   2484,11758,5832,13020,8272,8320,5704,6043,893,9327,6714,472,2788,6267,14134,
                   13506,10459,12549,1473,12401,6949,4613,11845,10001,15914,15634,9815,7698,3949,10336,
                   1757,457,3943,211,16004,12980,10048,5146,12228,12496,426,14373,13430,10312,10584,
                   5693,4293,3030,12300,3890,12520,12038,9493,5544,6152,7965,6297,7959,14297,8224,
                   11187,3779,4071,11679,13193,11295,8828,3157,12510,8434,12360,43,15776,10238,11319,
                   8023,4039,11227,16094,16104,5865,3272,12955,16049,8070,1036,4208,7807,4296,11516,
                   15853,14585,4031,5629,11971,11547,7405,3134,12864,14922,6144,13995,10132,9723,10701,
                   3385,2299,4372,5977,5655,15731,7159,4246,16175,400,1045,4135,13167,3621,8949,
                   9696,15233,6631,16103,13655,6733,12263,4003,10020,15418,3425,5469,5970,14461,6730,
                   3064,12905,743,15674,2469,1863,2605,10374,2700,1383,1827,9590,3435,9782,8926,
                   10248,15101,2663,11707,13503,10741,3011,10816,7247,9232,7357,11497,15269,5687,2471,
                   3968,4475,13606,5243,4004,14025,4111,15709,14417,9534,14930,12127,9797,12006,13205,
                   11697,12205,14914,15829,4588,2300,14980,2004,3319,15108,13791,4214,966,8461,10882,
                   4585,4200,14781,13706,13078,4226,8968,4512,8156,8479,2945,6275,3937,14200,2563,
                   3790,7054,3367,14366,9905,13296,11834,2539,13619,8246,3439,11504,10088,9505,10382,
                   961,13351,9482,11347,10058,4314,7056,5764,16086,1338,3699,1832,14963,14998,6195,
                   6107,12023,3559,686,10377,7022,14146,7816,9293,1327,13391,4172,6985,10509,9761,
                   6172,6137,8513,4424,5723,14121,11493,14758,8352,15165,9889,15314,6253,12235,758,
                   9538,9587,15502,7910,1925,8840,14727,6541,2649,8143,11013,15065,12849,3934,3744,
                   8883,15973,14849,12299,3487,10297,15590,12736,1897,15316,9471,201,10823,13820,15464,
                   2614,2258,5858,14782,1648,5064,14437,449,15385,5944,14616,14487,12807,14691,8996,
                   931,6500,2380,5211,2843,7688,11129,8951,13285,14911,12916,4514,13657,1688,7393,
                   15827,13437,13751,12028,8707,12975,9651,11659,9393,3880,14292,5005,14842,3576,11714,
                   7746,10410,11047,11665,4059,15234,13168,13803,5405,7004,10616,6916,9220,15349,2817,
                   10427,1911,5830,5841,3719,11213,14615,16085,8302,15288,9,1115,16378,8943,4531,
                   8131,12362,485,14465,14357,3799,3504,5362,14843,4962,9435,11350,3899,12539,9498,
                   5104,16271,14313,7145,7131,12057,8041,574,3930,7487,15713,13326,3600,9314,5505,
                   2158,15032,9076,9700,447,12085,1104,4487,8373,12957,10994,15718,13961,3853,6764,
                   8367,13045,10641,9686,6872,12537,9915,3069,12347,15762,13615,4107,4320,13860,508,
                   7668,6280,11874,6591,12010,13577,12237,10031,4926,14436,9446,81,10246,5728,15883,
                   1271,175,1502,13913,2829,6809,7059,2419,9122,11683,2493,16322,7307,5603,325,
                   13377,14188,3815,9111,1088,1333,3737,3313,1646,9133,15479,5154,8098,6299,5307,
                   1095,3637,1914,5011,9499,1605,11755,16047,2349,6971,15694,10853,3181,13474,1455,
                   870,5347,8522,9388,7262,8174,2222,10136,9542,1133,2415,7875,576,15309,15082,
                   15171,8259,14997,3735,756,5862,16207,8649,3024,12096,8739,14226,6552,15645,15655,
                   4658,12229,6972,2016,638,1638,13312,7269,5097,15478,9328,11402,11608,7769,2999,
                   4245,11344,9901,14020,13368,15684,14528,9300,11190,2672,1743,2960,3154,14532,504,
                   5928,4442,5601,8894,4597,1693,3059,9144,15079,11774,12827,9526,1374,10557,15962,
                   9690,8710,11332,8647,8202,74,10513,14420,2534,12240,13134,2094,11120,14988,9934,
                   4439,12842,13922,13603,2381,4939,1137,5632,13018,5792,3432,11595,11338,144,1420,
                   15379,10510,15810,2867,407,13283,11419,11197,11717,15381,8128,1496,6820,5908,6400,
                   14799,6227,6033,15764,702,8229,13607,4789,6869,12603,450,189,1906,878,15397,
                   2325,4503,6824,2051,10444,150,1686,9711,668,15513,9463,13518,4259,15292,9017,
                   10567,740,14875,3499,12020,8501,9104,475,5374,3633,558,3715,2750,126,12569,
                   7640,11579,1482,12612,1842,2928,9847,9036,12797,6201,13897,9330,6390,13624,10894,
                   3270,13817,11184,14156,6620,96,6564,12950,12082,11950,1094,5100,9952,10746,15529,
                   2286,7987,294,1161,3328,4403,11598,7834,13352,8619,15034,4381,14283,7550,3164,
                   11123,11580,12833,13965,11387,2332,5608,1587,438,10499,15898,13355,15986,2902,14855,
                   15190,12719,13479,2585,3306,871,5117,12410,14807,4023,14100,5549,1834,13477,2836,
                   7845,16022,12637,15002,6790,11961,5003,3505,809,1679,3091,3342,1493,8614,6020,
                   3921,11380,10618,5274,3632,11565,14686,12163,3060,14704,8109,8556,12018,10847,2784,
                   9473,8234,12659,3868,11964,2780,1416,1082,2739,3747,761,11520,8134,11154,2382,
                   3655,691,5445,7005,4974,16011,11947,9556,12814,14349,12217,12110,8354,5546,7256,
                   4436,11367,7712,12642,534,15173,859,5570,153,4482,6360,12845,11661,11163,15782,
                   1408,5759,9421,15145,11927,6687,1544,3167,1448,11700,9630,239,8105,690,5403,
                   6375,10590,3730,12137,12369,7574,4549,1302,3727,11116,10950,11169,8907,9078,6170,
                   1621,13443,14718,12811,15162,367,11703,5971,4752,11276,11095,2169,13378,13171,10912,
                   1873,9811,2697,2833,7092,1976,15115,6497,3429,6947,540,10787,608,2791,7985,
                   8755,16006,5715,9445,14709,1297,10072,7291,3605,2639,1117,8734,8280,9315,5025,
                   16284,374,3557,14426,14269,1705,1411,15217,13194,1477,5846,9196,14601,1600,8329,
                   1711,15626,8035,7523,11435,4125,5892,12690,4570,7028,14037,14230,7453,1879,3941,
                   9677,9941,7097,8846,6893,707,9807,15160,4674,6153,5414,7257,1835,5352,9885,
                   14236,14484,9183,14106,13700,11627,14381,10910,7518,10406,7737,13695,8785,431,6113,
                   7294,13086,10405,1046,5423,858,715,15241,138,6722,11053,10798,8909,10547,8977,
                   8027,10393,36,4557,7673,4098,355,10845,9101,7566,7700,10596,1025,13649,10338,
                   9109,6965,8139,11601,8895,5178,324,5084,11316,1550,13935,4469,5332,1586,9775,
                   7656,16170,14845,5820,6710,655,11969,6027,14814,2947,11055,15720,14400,9765,13394,
                   1713,15412,11970,4714,6265,2032,5213,1136,2490,3823,7801,13665,10940,15359,3804,
                   15804,11610,6977,1378,7962,4523,185,8572,1633,803,8086,11733,13811,15730,4730,
                   6956,12231,11208,3005,11949,14578,6393,15228,1348,3045,10386,2276,4126,10436,14570,
                   4454,10324,3669,6738,10014,6089,8322,3066,12477,1305,13729,2863,8874,11557,4340,
                   2470,4784,4086,10243,10744,8334,4292,4666,14149,8766,4500,8660,8030,9213,3175,
                   10314,3388,8954,4627,8321,2185,15416,15031,9095,6319,12660,1905,1012,16007,5493,
                   7850,15044,13513,1706,8345,2437,14120,4880,13172,15552,2841,2611,5069,10247,14636,
                   8708,203,6713,2612,9092,13541,9917,7665,6251,4156,15060,6576,167,133,4104,
                   14093,15383,13067,3461,15665,6189,9684,1006,11886,12050,14153,197,9420,5432,10794,
                   4206,11299,8464,4853,7057,8607,15951,15119,512,12000,2796,4358,14808,785,3539,
                   15568,15202,8682,1655,15792,2290,14077,24,5946,7546,3393,1641,12667,2966,10654,
                   11908,5215,13019,9257,10733,8502,6866,14060,10634,16276,7696,15236,9008,10316,11284,
                   15640,1275,15679,12195,3146,2488,13609,13339,7265,10335,7224,5950,10193,15387,5614,
                   6711,11852,8218,8998,15389,12270,16247,13189,3363,4983,1910,4623,11759,7990,6750,
                   13114,2633,9517,9043,3718,4984,12171,3153,14881,3419,5516,9197,9067,7676,10880,
                   732,5955,11583,15283,6285,2643,9930,4923,2259,15823,963,5136,16206,16105,4701,
                   12199,13631,9143,15081,716,16035,6349,13829,8587,11069,7997,3208,3913,9244,9771,
                   16318,1539,3406,14174,3187,10807,10370,3137,8532,2413,16313,5527,4124,2810,16018,
                   13765,9779,7663,6670,515,13709,3115,583,7666,1038,12396,1402,5234,6401,6480,
                   4252,6547,6476,9218,8780,4019,9674,3381,6992,2586,13770,9224,11687,140,15546,
                   11644,7194,5176,4443,16377,11709,10607,6474,6333,8436,3887,10116,3905,8081,1762,
                   13111,3055,11508,4930,14617,5784,7547,14029,14027,5817,7225,9019,14163,11582,5852,
                   3522,15516,7380,8808,15255,9477,15893,12819,3594,15663,6165,832,6521,8590,4753,
                   5468,1342,14679,13733,10610,4373,4729,7456,9607,13582,7226,10780,3338,1308,11256,
                   13621,6522,13720,12674,4476,11407,3168,3679,13636,14198,2122,9467,2580,7394,11540,
                   7026,7718,9598,6179,10120,14104,791,14277,10766,10540,7116,8714,13667,9908,2895,
                   556,15284,11573,9344,5370,3920,11125,14495,9139,11510,14815,5618,16080,13772,11995,
                   12381,15765,5238,11737,13307,7680,13804,136,4275,8692,10608,892,4628,9023,7863,
                   6462,8546,10280,15068,4324,12868,3162,2040,14954,10824,4290,2388,2225,1505,2334,
                   7781,14887,12517,12626,12902,8173,2845,7462,12625,4573,10367,3104,433,11001,9991,
                   15450,3680,7661,908,15897,6122,10127,12727,9185,6304,11559,8475,8323,5676,10545,
                   4553,15570,1677,12725,14286,7652,15935,3497,11839,11997,1291,12485,8037,4599,11035,
                   6194,4861,13403,806,2971,3525,430,5565,9318,13914,13309,12504,2591,9195,10400,
                   14078,6081,15896,16021,3507,10785,709,2378,1487,6452,13464,2839,12179,6238,11652,
                   6173,4877,2524,16230,9415,2105,13278,11399,4721,14923,13396,9565,12281,12355,9338,
                   8994,4675,5545,910,3099,10143,8283,1034,9087,434,10233,6662,10045,833,5966,
                   1040,13681,14560,15,5460,1620,4876,6136,713,1063,13950,7091,10121,6004,9382,
                   9994,2683,1619,15150,320,12900,11041,15664,5751,6647,2195,11341,7284,6106,4860,
                   9190,15321,11812,11091,13896,5290,13140,12412,14396,10696,12406,1748,3036,4528,216,
                   12321,15753,7933,59,2133,7234,13863,4128,12650,2099,7304,9085,15583,993,3722,
                   14798,5237,291,13317,2951,1031,1801,10047,9054,8351,7326,1197,6134,11653,14392,
                   1453,16072,15936,15325,12071,13737,6300,9320,13727,7664,5739,12234,4888,3475,9378,
                   13061,6447,12303,4496,9342,6606,8120,15954,2033,5630,14135,4634,2359,7796,15105,
                   4481,12939,974,2944,4827,4567,3295,15337,2529,5057,7669,15266,12513,15282,5855,
                   10215,13525,8471,794,3837,9113,2905,15932,9981,7645,7964,4677,8099,5099,6247,
                   13736,4074,2877,6085,9184,10568,9969,10299,1009,10217,15735,14926,12128,2344,1446,
                   7238,285,12661,5710,15706,10838,3742,16002,3026,12438,8669,7330,10311,7738,11422,
                   13983,8437,5934,2719,13375,2996,11978,1839,8359,3784,8775,1195,12115,13899,11056,
                   16329,2306,13828,5872,2850,6777,14507,6831,6682,35,220,6385,15623,11535,5426,
                   12844,11229,2911,15976,7254,3364,9511,9826,14272,918,1294,14734,6826,10591,5446,
                   825,9851,65,15567,7809,4041,8983,14430,221,6357,978,6987,11945,670,5293,
                   9331,15229,5662,15530,13598,22,1495,729,2109,5235,5909,461,13679,3650,12853,
                   9335,10818,7613,14443,1376,14229,10831,3629,1256,1367,10587,3194,3998,9070,9949,
                   10414,12722,8005,12787,2830,7302,15960,9103,13752,10201,10365,9438,4229,12102,14196,
                   16337,8018,1562,14255,9049,15705,10897,1864,3553,4045,13060,6257,7011,10329,12372,
                   12130,6130,13465,7836,9519,13754,10063,9892,2695,13380,2196,6046,8547,4545,14000,
                   6706,6622,3961,1950,1289,7364,8383,14062,5933,10606,5913,6546,1323,1463,5910,
                   4253,8750,8529,13924,9731,7007,3879,11363,14576,9312,1845,15983,12047,7040,2202,
                   15114,5483,9203,8181,4937,930,4202,14960,4222,694,6616,15540,3544,10428,9248,
                   7572,7322,8265,8075,8611,7924,3489,13015,7771,8591,5968,5987,13620,15769,115,
                   1565,208,15214,10071,12892,2885,14005,6920,15799,9469,15110,14353,16090,9640,2648,
                   4898,6908,11134,2351,14738,6477,5912,14858,6788,7128,2530,5143,14227,9665,3526,
                   4495,11672,7248,4565,848,1237,4363,16064,5302,12951,16219,10402,11593,4250,12404,
                   2635,12391,2431,13556,1779,5742,166,14320,10915,786,13348,13459,7240,9944,4353,
                   11448,2477,2283,14499,11875,5059,14334,10457,6724,327,8063,11028,12531,2814,797,
                   8733,7971,15996,4400,942,6261,9343,16225,7373,7165,3430,10321,10235,1292,11841,
                   6506,15541,1856,1119,5300,97,6467,6707,1868,16305,11219,792,4133,14647,15232,
                   4743,13522,9125,7135,3409,8651,15106,11077,12284,7505,7543,12351,8243,14818,3015,
                   2194,6190,9672,3050,14731,645,6755,8179,9713,9497,10304,589,580,15444,3975,
                   7150,6162,10044,8483,4327,8517,14407,12601,11795,5899,7662,14203,7929,13162,1920,
                   10638,14453,14127,3451,7755,14311,6354,34,10330,3359,1545,5436,10905,10946,12920,
                   2173,11321,13686,2189,2652,3978,11250,12292,223,7636,1614,1972,1157,7716,7103,
                   6466,6623,14018,7410,5615,5821,202,5733,4631,9326,13836,12899,12079,10873,1938,
                   14013,5575,139,6594,326,10563,3821,3183,14482,4755,14460,12262,4746,11089,2336,
                   3590,10228,5674,10015,13806,6988,3571,980,13843,7003,8381,14828,4405,11919,5835,
                   7991,14308,9272,8178,6652,3414,13590,2013,10524,12169,13264,2959,8039,5040,8366,
                   14692,10077,1149,2508,2363,4020,13886,298,409,3443,2851,6351,13148,6822,15265,
                   4399,3803,16166,820,16134,2893,11893,6549,14859,5360,11960,8891,15998,11305,13514,
                   8072,2280,7482,12790,15149,10373,14754,9576,11383,4166,693,16229,7058,5076,13046,
                   14150,10588,15166,769,6927,3567,7536,11988,776,5233,1497,6779,13149,5253,4502,
                   6373,14735,3378,4027,14506,6353,15600,85,8468,11575,7440,4271,10571,920,2082,
                   13611,4159,13386,13909,14891,15682,227,15420,4369,11110,2570,10079,9638,1028,3767,
                   3473,771,2742,1081,11976,14747,3582,3217,2608,7382,5797,8503,12602,5244,2384,
                   510,5045,9687,7777,11451,12858,12912,11093,2706,382,7207,2087,9745,204,11842,
                   12058,597,4225,3695,12755,12573,706,5540,15816,12873,4171,14066,7947,8294,7063,
                   8865,12074,13480,7815,8171,1777,8089,6542,11135,9838,16136,16191,9891,12696,1913,
                   4977,10617,13432,7839,6533,14004,10523,12379,14736,2933,768,6815,7335,7623,10108,
                   14470,15697,15207,3677,4178,9064,2401,20,16128,12575,14410,9939,13544,385,13853,
                   3428,5485,12400,4641,3127,7126,7961,3692,12311,9261,5656,12230,7329,14222,8286,
                   10416,12968,7174,9108,5597,14878,8936,12717,15523,15695,5110,5148,2017,2455,12352,
                   11611,5643,11931,15543,7704,2689,8195,10203,4173,4873,979,6387,6741,13807,14674,
                   7549,5919,3380,3049,15305,7437,2921,10347,1576,12930,13333,13842,6745,4975,5404,
                   3878,6486,2501,13416,10328,6448,8010,10715,10711,1419,16067,14314,14058,14717,16320,
                   16365,4866,14147,14633,13489,6001,11541,5530,14036,11596,12946,2150,13794,1229,16220,
                   14361,1685,50,12242,6494,2203,4130,8307,2978,14761,15471,4195,1485,15549,10702,
                   1613,12012,11108,4832,3366,4852,5765,6808,5077,11444,3762,8864,6900,4607,16063,
                   1535,9270,997,8123,526,2913,8934,9734,61,13622,392,13161,10598,14322,3788,
                   567,8100,631,14681,8341,537,11768,3254,3074,13951,6177,5480,1977,10174,12607,
                   8847,5538,12870,11990,9658,15856,7717,6705,2022,7728,3222,8778,9375,4415,15526,
                   13918,15884,10284,2754,11064,6011,10541,11102,12215,2061,1474,12489,16334,3782,11181,
                   6951,3126,6550,2531,7144,5015,11417,16251,3408,6634,12738,15238,4189,2600,9163,
                   8760,3371,12190,7130,5014,9922,14017,15916,14073,6661,3974,2482,15493,13504,15508,
                   15199,14034,4247,4732,13156,14158,1057,14777,3431,6610,1608,13184,8672,8852,1211,
                   2143,4118,2881,6963,12969,12877,780,7596,4568,3368,11349,12763,9668,308,3397,
                   11437,14404,2982,12331,7831,7276,15991,4095,5927,11645,12480,13109,12408,9919,11246,
                   16000,14374,1739,1558,13882,383,6881,3645,8486,10396,2802,16130,11018,15860,12766,
                   4379,3346,10130,14490,8859,15224,10997,11293,5816,5951,5981,13583,14630,8326,13462,
                   3807,968,13441,6216,13862,14978,3687,6316,284,6583,13458,11104,8271,15650,14438,
                   10817,4779,6558,4564,491,13487,665,13660,6365,15977,5415,5547,11943,2735,4063,
                   240,5120,8175,10334,5814,10348,951,13313,5153,9072,3951,8604,13831,2551,10615,
                   7191,7830,10757,13793,12336,15147,10805,9081,6193,11340,2156,9703,12978,11322,3604,
                   5498,8060,2343,5566,13087,2174,1107,10083,12919,3202,3244,6426,15961,6221,2098,
                   16323,5083,9862,10421,10413,10891,4146,13799,14051,14456,11555,7600,11460,1085,10909,
                   9575,6512,8264,1858,11681,6236,1196,14223,6958,6327,8668,8637,15774,7622,6928,
                   13835,13980,10549,2686,1387,3402,1212,10754,12333,521,13532,1073,8192,2665,15561,
                   9903,10760,4310,3467,16096,9233,4781,10645,10926,10751,1817,15372,337,6471,1288,
                   11637,12744,13848,13090,1110,10245,16224,6609,11267,569,14889,13604,14241,9766,5958,
                   8809,6865,2609,12213,3096,3980,11291,2112,9643,12117,9848,15826,4950,5999,2581,
                   8629,11097,2428,12452,4042,11303,14285,9397,11546,4717,9925,11238,949,13288,6709,
                   14019,8743,12339,13494,10753,4526,12469,14133,8415,2297,9926,14869,16158,9303,8526,
                   15179,13037,9014,13096,10351,253,1831,8947,14973,7857,2920,6996,11165,13932,6836,
                   4270,2295,9611,11785,10475,496,3761,617,3593,13335,15875,14231,5533,2727,9099,
                   5978,9606,8056,15127,2724,9440,6068,12624,14895,9592,258,3530,9051,3780,2567,
                   1220,1656,1238,2546,3293,4076,12108,9173,3888,13006,12653,6798,12791,3161,16118,
                   15712,5020,11189,14472,9614,1125,1369,8677,10408,2165,15559,11721,1223,9718,4211,
                   10718,7731,15310,7542,6640,9561,4617,12783,12313,15539,10291,985,4384,9193,847,
                   10054,10642,5559,10911,8921,625,11434,5524,12267,13801,13435,15121,15667,4298,11482,
                   12563,8227,12463,12098,3854,6817,3566,8792,8125,815,10260,7504,6641,14751,9020,
                   5785,5947,14675,6991,5324,3165,8960,13274,9620,13072,2035,12992,2341,1026,11447,
                   2441,4525,16114,3562,13903,5590,7701,3170,2391,4387,7634,6511,9249,5451,12368,
                   3540,16201,283,15485,11086,10930,1281,13626,15812,12693,1070,2421,9965,8603,7879,
                   8922,926,1527,8748,10682,7178,4569,11237,10725,7317,11554,9795,16099,15794,8919,
                   3391,13056,2820,7926,15615,2355,14442,6408,11326,1358,13260,9942,11604,14274,1428,
                   16106,7334,6929,1312,542,7684,3659,4555,13929,2544,2177,8796,12564,7571,4386,
                   6700,1615,1352,13759,5281,12568,12034,653,9980,6295,10528,2273,16215,2121,9589,
                   15880,6096,15934,1154,15006,5611,9774,9830,13389,909,6078,6671,5898,6250,5738,
                   5904,1039,5056,6281,15908,3765,4556,5585,3145,1644,5849,9066,7916,4409,6036,
                   13805,15576,3892,7626,3658,14724,11513,4941,2842,16258,10843,896,3043,525,4237,
                   5801,16277,4648,3948,5591,7567,7855,8221,6980,2688,11254,16014,11414,9500,13696,
                   6,5418,12643,7846,10223,6704,7102,6002,9599,1113,3009,13318,12385,171,12152,
                   12577,12971,7105,2023,15311,7502,9840,2641,1121,8388,10407,5561,6329,10310,12571,
                   10575,564,2977,904,380,4966,10411,16149,4304,8666,9786,1680,9034,14310,6680,
                   3503,9951,11914,2116,2480,10011,14795,14220,4574,12788,15049,13781,11609,5159,13014,
                   6519,12771,11850,2968,7811,11450,6874,4586,8147,2335,6061,14933,128,11552,12184,
                   15437,3000,15364,8520,1775,699,14505,9068,15263,9824,6269,2358,2504,3702,13664,
                   5636,16101,13301,990,8795,4297,4708,4040,6380,2969,7775,15015,11044,8170,6904,
                   4868,9292,4092,8499,11612,13347,15887,622,12335,14488,2939,15995,4478,2778,7277,
                   7190,12376,8598,5318,13353,6454,9518,13433,6919,10723,13692,10332,1806,16023,5356,
                   7714,10222,12943,3683,5716,15045,755,12640,8220,7702,14972,7435,4155,10074,11244,
                   16083,9022,6045,8191,11308,281,2963,2452,292,9585,10791,14749,13345,2414,5127,
                   15864,13251,8923,7590,939,10100,10478,14907,228,8015,11063,14666,9386,3284,16373,
                   10860,289,10257,9537,9365,11560,15208,11061,3515,13209,2201,11282,10307,13931,10446,
                   15168,4069,13788,12297,4894,1924,2180,14784,9178,3809,7678,4408,4456,2252,8686,
                   3884,3234,2579,6516,3488,7609,2821,14202,6673,14428,3910,15752,6213,13921,4142,
                   2393,11375,2237,8576,15302,2540,14224,1246,778,14409,8295,6898,12246,10672,3330,
                   12325,235,9117,15340,15801,3348,9290,14296,4678,3693,6952,5645,1379,6296,4676,
                   12586,15306,12486,11073,15997,6602,16138,15565,882,1919,8530,12526,479,2720,12854,
                   10380,8433,183,8754,5490,295,5312,12728,2387,5834,6751,8887,10676,9987,8188,
                   3209,5876,13206,13586,14402,12646,9310,10984,12723,6423,2374,15414,2395,11790,7012,
                   10714,15043,8984,229,7885,1202,1434,6437,16336,8476,2479,4038,4696,16142,2714,
                   8976,5581,4072,9175,5698,9212,13126,11157,15627,5523,12484,6103,2958,6763,12056,
                   5017,1181,9708,14763,13076,2675,9398,14710,2247,9131,12015,9400,15242,12151,12707,
                   7458,15126,14835,14970,7292,2342,11029,6596,13878,14424,9287,13570,13822,15944,4705,
                   16048,6796,2281,8610,6514,4011,1658,11021,14846,3904,5939,11863,13566,3700,11224,
                   5651,802,1776,6907,11959,12515,13501,10565,16239,2311,14707,2154,5098,6298,7082,
                   630,1662,11726,238,5443,8653,4240,14705,5381,14070,8562,14744,268,1384,12278,
                   16352,9485,2485,4620,6262,15955,996,7069,8793,7539,3630,10241,5231,15380,12363,
                   4996,1566,9437,5398,11155,16257,10263,11600,5598,1889,1159,11012,4900,4014,11397,
                   4587,7779,3151,12495,1438,4576,3738,1000,13703,1284,4824,8478,1261,11762,14040,
                   10164,2153,15499,4614,4282,16157,14246,16038,2826,7814,6905,2844,6066,5121,7263,
                   16232,3017,6754,6653,9202,6499,15297,15755,3909,9737,4249,179,7995,9986,11309,
                   7864,7348,2664,10202,6982,2793,9115,177,8511,14594,8972,5195,8646,9984,15440,
                   13238,11002,10521,15468,66,14982,10833,2219,2526,10250,8965,10424,5823,11853,7854,
                   7703,2396,13536,4680,11186,12462,7532,703,5241,15334,8418,4294,11939,5387,9472,
                   3586,13927,1440,3990,4192,14324,12350,6643,1780,15129,4840,3438,10659,14694,2763,
                   15047,2834,13718,13891,14638,3109,14469,14996,5132,3521,12989,4153,14068,7323,6513,
                   3314,13122,522,11139,11105,7243,4625,13021,9533,8625,735,2732,2270,16316,5503,
                   8735,10142,6157,11614,12427,6960,10417,12669,10095,16282,13406,3656,10628,6899,7946,
                   14775,13357,10889,344,15767,16189,4989,16084,14683,1700,4131,7043,12684,2593,3929,
                   12474,2870,13153,16203,314,14340,1546,3421,4165,4626,5705,5677,6088,4272,12095,
                   7229,14631,1710,5520,12830,3093,12139,14984,5691,10745,15926,11115,9530,10205,14680,
                   7085,3448,15895,2436,5720,3492,1959,9369,13551,9055,6235,4884,15164,5413,12111,
                   12202,12940,1838,6339,592,10992,9096,2473,2215,11360,6765,5041,14593,1086,4464,
                   3345,12956,5034,9740,549,10037,286,3569,10182,14829,6746,14063,6472,4120,9278,
                   14811,11030,7735,1120,12258,14096,13331,10835,12794,10736,1555,13642,348,3549,11081,
                   12118,2292,15557,3251,9875,16153,9717,15193,3588,15186,9127,10593,1634,14132,7419,
                   11024,16141,8231,15335,14030,2166,3750,15463,2161,10107,554,14741,2406,1624,9154,
                   466,182,7982,4690,12361,5935,6332,10230,12482,90,1442,12958,3265,3252,13233,
                   9082,13613,1847,13907,3444,10212,11083,9025,15274,14102,12366,16267,11953,10922,10883,
                   4814,12545,15205,5763,11298,1278,3481,6834,11574,795,6288,262,14141,11558,6087,
                   8020,2478,8157,4825,11764,10887,4326,6664,13385,13372,7209,3644,1499,12673,10293,
                   2328,11039,801,3579,13052,89,1598,4093,7819,12021,5271,5796,6867,10666,12803,
                   11913,1760,14541,4537,176,8199,4425,4878,4466,14145,14406,6666,10342,3500,7789,
                   15365,5118,9389,9161,13973,7425,9302,8751,6483,7976,12527,5889,3136,15580,9158,
                   13150,13812,12679,12915,11433,3924,12155,1841,4162,14459,6047,6463,8805,13447,10730,
                   12186,10879,725,302,14074,5382,12019,193,10362,12421,109,8111,14071,11731,11022,
                   11042,9285,8975,11252,2138,4186,5648,1632,181,4221,7939,2236,9522,9479,3028,
                   4451,9867,15139,2846,10952,11068,5874,4116,10775,5969,6520,11027,16280,3903,1981,
                   11413,9828,7833,12377,1758,11424,9964,7589,7272,13830,15950,5766,11523,2102,8074,
                   6515,9689,12464,5369,1492,13529,2521,15035,5320,11389,14722,14117,3405,9532,8275,
                   14864,15447,11096,7396,12676,4364,9929,1789,1603,12982,15775,7332,907,52,11263,
                   1017,2053,11491,2106,9625,8203,5194,3025,5138,15107,6636,4241,8106,12069,13516,
                   14619,13946,15458,14307,5697,4501,964,8905,15112,12528,7750,9787,7331,6326,13597,
                   3740,7168,8853,12799,9790,1368,7493,4434,8844,10555,9569,5778,1654,15849,3259,
                   7920,3885,16303,2289,1397,886,6040,10609,2275,2607,1824,12809,1346,2312,9013,
                   14186,12681,1893,12621,12756,12029,4955,5731,14637,5192,11333,8839,10134,6012,13666,
                   2886,1571,16077,1478,1978,13242,507,11427,15681,14033,3281,1697,13050,14793,15075,
                   1782,796,6601,5502,8281,15423,2,12097,5141,10163,9982,12338,7412,2364,11311,
                   2988,14913,7594,10683,6482,8528,12710,2254,7984,5491,9384,1316,3608,2918,7141,
                   9162,2661,1812,12428,15013,5695,14148,11405,1695,492,11514,11464,9834,3785,6341,
                   9308,3128,7107,3223,5915,9219,13398,12768,13694,5563,834,16028,15904,2874,10884,
                   1730,7538,8124,991,7805,7632,12565,12063,14862,3302,12523,9206,11488,13446,8548,
                   2658,15669,5959,7381,3374,11671,13777,10848,594,2410,11607,4505,11486,662,15448,
                   169,10144,9961,16374,1103,15966,1727,4687,11294,12227,10494,629,12829,13190,10170,
                   330,164,10135,8712,4896,14726,2115,3580,8679,4435,5539,7096,11174,12275,4256,
                   8933,7169,8673,10932,3337,14377,1490,15225,7220,2091,2369,14412,1810,7062,6901,
                   10811,2486,4339,2737,13159,14193,2708,15425,5683,2862,15156,15732,2603,12634,12456,
                   15784,15972,4906,10301,318,10677,7992,10017,9661,15999,6792,15063,15017,5179,5600,
                   376,9856,9323,212,10187,9304,13027,12804,965,8663,9079,5458,10546,5578,15956,
                   4016,3959,15357,9799,9996,14500,10123,15795,7605,624,7520,7591,7878,103,13769,
                   4770,10249,4185,13888,1672,14435,4257,8851,7072,9735,6967,14879,10450,3101,8989,
                   13548,4530,4994,15185,462,1830,7433,9697,4740,11128,4943,2995,12146,5703,3389,
                   3914,14555,10060,4268,7552,13275,11806,15593,10425,8216,76,13314,4822,4513,4604,
                   13774,8201,14595,11253,8568,8026,5580,14673,14629,12423,14896,14431,6382,8013,15042,
                   14166,323,13549,8940,3278,14497,11800,12895,6151,9339,4935,14690,5824,15388,2848,
                   16061,13003,464,12149,14172,2626,4103,5803,15237,13081,1325,14187,8700,7428,13097,
                   15293,5265,14162,5952,7545,14750,7862,6044,11082,8453,13221,12254,11144,12348,15131,
                   14599,9967,2914,7753,1681,5288,12796,1259,4417,186,11015,9516,5839,92,738,
                   2823,2757,15704,6440,3781,7468,3708,10792,6234,8350,11777,9216,10191,13302,4471,
                   632,11232,15286,6936,2400,7677,5848,7793,14504,6419,3999,7270,3950,12991,1100,
                   5028,9701,5459,8906,10804,7283,8446,13612,15582,6222,1035,6159,14713,12328,3232,
                   13413,5735,2613,15030,5709,8362,2472,2726,7455,10844,5589,13753,6428,5272,474,
                   10692,11353,6964,5596,3814,5089,3836,6291,2792,8197,234,7953,1364,9258,13714,
                   13628,5079,2418,13523,6633,15187,8411,11273,11548,12014,8050,1647,5095,3138,13200,
                   11300,1561,11511,6024,10477,10728,15080,5868,5183,3058,3035,14925,3882,12752,15067,
                   14967,11722,9692,8430,467,15181,11587,8535,15581,13972,8524,8761,7140,15453,15024,
                   247,198,10773,12448,2408,14136,3889,7478,4073,8029,11075,12618,7914,3808,9573,
                   1985,14485,5553,6305,6084,16079,12053,1855,762,6196,15320,846,7514,2590,6119,
                   5517,5847,3052,12389,9872,13875,8180,6498,15760,13217,8802,11489,4485,9645,14534,
                   14816,8031,5699,3532,3071,9057,11776,5914,8781,4978,15348,16296,15055,5922,11686,
                   2321,9376,4082,14968,10876,15102,4780,7356,11400,13281,14553,11307,13456,10226,11770,
                   3672,1242,260,5879,3912,2916,15981,6510,7573,4136,3640,4160,11355,2852,4371,
                   10732,5794,9119,1365,12310,6955,3357,405,236,864,1394,1219,11804,11261,7067,
                   1534,6753,14309,13900,13187,15011,3321,8385,4121,14873,1461,12211,14253,11043,8567,
                   13571,8066,12713,111,7957,3349,7817,4869,12554,14950,3849,11603,9623,14543,5168,
                   11191,8527,7424,8901,10186,9618,11071,8776,3129,8002,10985,6490,1844,5024,5504,
                   2573,15992,6114,13915,6248,13726,213,8898,15923,3477,6715,4630,5156,11403,5292,
                   6391,10559,62,10819,6406,1515,1866,6150,8995,1945,14959,6260,6607,6019,11572,
                   12459,14370,2772,10829,3076,1821,11695,13270,11885,10199,11690,3286,14797,1215,4112,
                   9502,14328,10968,9536,7895,9682,15815,13550,8348,15333,2953,13358,14447,4414,7108,
                   9227,2320,6255,3474,4217,365,6180,9995,8756,1317,7888,3285,5119,8523,13370,
                   3103,11658,4959,9666,3599,14284,7403,8047,2674,8052,15243,10581,11836,1636,9452,
                   15212,437,15737,1227,4035,12222,518,11811,2104,6140,11550,244,2148,15059,5758,
                   5433,15575,1501,15965,12888,9726,11016,10463,4065,13632,11235,13484,1335,11351,5006,
                   1567,8133,6432,4228,7461,2725,3072,11498,14708,5494,5066,80,12508,13712,14023,
                   3225,9405,1637,9820,14841,2186,13034,10637,3916,10538,12196,15512,5261,12250,10726,
                   2123,5997,15798,6535,200,4916,8235,5386,10802,13257,15254,5961,9523,8579,13147,
                   9887,4848,11346,16353,8117,11986,13868,15698,15605,14474,4440,12039,4673,13778,15920,
                   9712,6655,5010,5105,7709,11415,9361,4113,10383,4844,2985,13043,15903,14898,3365,
                   6367,1532,11357,15125,10998,9042,5838,7837,6455,9971,9571,8578,9478,10039,1964,
                   5187,12826,1350,10550,8338,10204,8624,8274,4795,14416,9364,7894,4891,759,4463,
                   207,5124,1132,16223,4280,10002,54,13564,4490,14462,16185,14043,15830,10176,15443,
                   5408,12815,11270,13454,4616,7506,11391,4382,13397,6147,16371,12580,10554,8681,9970,
                   9521,1984,9180,10908,7321,6803,14755,10268,1032,2002,10184,14661,11899,10790,7870,
                   15503,4892,15881,7650,4767,1826,7465,14894,13710,15342,12547,486,6003,7719,15339,
                   11876,13561,16368,13815,11756,7457,5979,15563,10742,2294,7443,1150,1199,7490,1124,
                   1002,9656,9306,11070,7554,13073,14542,9298,2107,8645,483,2030,12967,12936,5441,
                   11701,10965,16293,2100,13005,16127,3299,6853,10078,6539,16091,2113,7389,4484,9209,
                   2256,9895,4078,2523,12974,4957,10209,11241,11872,1949,9617,1003,7100,15857,10016,
                   8889,1895,14161,3527,6554,9394,3598,7183,12762,12665,12890,6648,3051,5917,4018,
                   9940,5536,14520,3984,4123,3561,9366,15814,5752,1007,5044,6873,12465,8612,5191,
                   15963,9153,11723,14386,1575,4741,8948,13320,2330,5029,9077,2157,7287,3528,13617,
                   2882,1916,8043,1180,669,5258,9496,6654,916,10707,16152,8407,7499,1222,11832,
                   14569,10700,4724,13658,1578,9426,11017,343,3863,13925,6485,3511,15298,7073,8935,
                   3908,8185,12295,12430,8374,548,14342,15319,2086,6883,12165,12775,13991,16324,12593,
                   3983,3086,1427,10717,14990,12929,10944,2212,13382,10508,4875,14773,1991,13395,5624,
                   7379,14240,4176,10827,16319,5880,12657,13827,7657,5610,11799,3334,13764,5897,379,
                   10271,4769,3434,12440,15741,7751,8667,3955,12282,8675,12798,4420,4231,16098,7602,
                   12007,4798,9997,8914,11718,2319,14243,736,16205,830,15161,5542,1967,15294,1872,
                   5477,13176,16146,15635,4647,16161,1953,14884,15819,9454,14840,13885,12617,7795,15262,
                   6368,14273,8597,11412,7658,13388,12382,13071,8773,11465,14082,15802,6910,16137,7732,
                   2640,1307,11469,1129,3870,2929,5287,7391,12116,824,6377,2532,3470,15891,15876,
                   8897,377,15405,11639,2972,11569,7308,10420,15978,1022,15138,8582,16016,15872,4498,
                   11649,9200,13874,3250,8405,1190,10801,10252,11780,10156,11453,3844,15174,14237,5550,
                   13146,9481,15315,4886,16190,6913,6458,2694,2257,9647,14477,3159,844,10502,11345,
                   5163,15560,7351,14367,4835,14586,15116,6014,2894,13088,10218,15222,4144,12536,5047,
                   13540,5737,12409,7199,1940,826,7146,14016,11239,7406,7421,2296,1788,8632,5857,
                   2642,3873,1809,5205,14989,14258,12558,13545,6942,9676,5537,7617,13261,6584,4352,
                   14548,15051,10415,6420,3502,7757,5308,10747,3458,11442,4610,15122,16347,3032,10145,
                   8823,13948,586,8602,7588,2915,9032,10569,6307,9570,9520,14279,1301,16042,13174,
                   15691,2679,4151,16236,7644,6294,8741,10162,8204,15441,8189,7994,13142,11674,11000,
                   6075,11712,15466,6181,9383,8915,9798,15969,4376,15915,4644,9546,55,1752,14698,
                   2681,13581,16092,3484,2481,7761,12364,2671,5675,6739,9660,8888,14940,10093,4749,
                   4002,2552,3211,15846,3047,14805,14790,12245,10688,12236,5063,13741,1193,11669,3994,
                   287,8376,1965,9524,11454,14766,15505,841,6663,6163,1800,6233,4657,12981,10465,
                   749,1079,14573,7516,10643,4538,10919,4850,4315,8958,4269,13755,6457,552,4351,
                   10978,946,12923,1099,15215,6529,5497,1296,7859,4154,14693,6767,9639,6852,3382,
                   13962,12918,7298,15195,10956,14057,2764,4843,11505,3436,15555,14941,10019,12668,8289,
                   10207,956,14908,3457,7881,938,14518,1468,10788,265,2160,8425,6930,14471,254,
                   13743,3834,14346,3140,13062,5937,3886,12030,13572,6005,6178,14501,8917,13767,12584,
                   12726,6082,2463,14142,7218,14491,4723,13994,8713,8838,5123,2223,2864,13850,15652,
                   3754,8282,6156,8822,9960,751,15854,14605,3212,10151,10150,12141,10958,12264,11531,
                   9880,11452,4561,12134,13552,14651,9983,8740,8161,14041,11364,4197,10448,10357,8835,
                   13191,14337,4337,7094,12606,9554,15442,13290,11193,544,16354,8379,3568,9581,2003,
                   9305,8900,823,15351,13303,9058,15386,5818,2577,11330,4049,13988,11884,9355,10364,
                   6430,8194,6983,9531,8339,957,10096,11240,9652,12460,13311,8451,3445,13524,6286,
                   15734,6310,9911,13089,12220,15620,7847,7715,14099,15486,9239,13457,6737,3591,8438,
                   12483,435,6161,10320,6613,4261,15579,4694,11318,3631,8127,4087,5689,1111,7371,
                   5068,5729,4771,8927,8215,2527,9878,11781,11584,11264,288,7893,16327,15461,7541,
                   814,16256,8137,12800,13640,16235,12454,9578,1033,378,9781,2931,16348,15750,2266,
                   12997,13273,1512,12649,6048,15069,13104,5,7113,15885,3276,4032,15535,14538,15538,
                   7511,2329,8490,13763,11315,3486,4911,1008,6308,319,8884,819,3386,6656,588,
                   11283,7903,11221,12599,7739,6328,4664,10585,5701,3174,5804,11285,11533,13039,10234,
                   6612,10859,14317,5672,3668,12663,14703,7010,6449,6684,3358,7842,1807,7264,5815,
                   4650,1756,5595,13648,1336,3372,8518,3501,1480,561,1577,6998,7266,950,252,
                   7430,2964,15280,2221,3684,10449,10169,4447,12780,10971,12209,8559,192,10200,6431,
                   4572,6071,16210,3967,5887,10806,15148,6801,4763,2604,687,4865,14015,3242,7981,
                   12855,4845,9504,4355,11463,5666,2277,12994,3952,4101,13894,37,5582,13993,11430,
                   7210,2803,1267,2234,6120,14079,6567,16218,1047,5568,5560,7736,7494,2164,4967,
                   7747,10890,7310,6421,9948,6961,8287,14512,1287,9863,7309,11140,13001,8217,8964,
                   2816,4981,6509,3545,2896,3088,1716,2092,13444,13137,5669,4127,72,16054,710,
                   15346,15400,857,5255,2050,7905,13930,10168,10356,8938,3100,15312,3172,13420,14265,
                   14335,6593,13507,4637,15403,11495,4064,9428,748,10050,3410,13559,2954,12961,3200,
                   923,16070,3422,11784,7445,10729,9140,7882,14906,351,2537,12851,1414,14514,12306,
                   11131,10704,12107,1021,15036,13337,225,15474,8831,12226,953,2027,439,5335,15411,
                   1345,9899,845,10986,2024,3412,12747,9760,4874,5222,15811,75,5197,843,13426,
                   12502,2361,334,12779,15469,8208,12378,6922,6759,2012,10864,394,7646,2272,13245,
                   11905,13954,16187,370,15924,16172,3266,9460,12197,6010,7117,12987,13735,4552,6090,
                   8908,5579,2687,7338,9529,1351,279,12033,9568,8680,1375,5189,63,9332,15021,
                   15481,3820,6726,13500,8093,741,5266,6306,9968,921,6838,1464,15352,12570,7741,
                   4518,2519,15071,1926,11837,9402,14597,12689,4665,10313,3195,6416,6812,15167,5447,
                   6374,1635,8412,14557,14114,5592,1024,7078,14323,3310,12935,48,4580,3282,15092,
                   6475,5932,6041,8693,5975,13732,547,15392,2550,7275,4976,6917,5373,11381,15477,
                   11900,1143,13422,11704,10981,147,15739,8293,3657,1664,15901,10936,1887,5799,14061,
                   3917,9458,6676,14452,13044,5043,7517,10055,10927,7358,14788,3509,3775,14052,1582,
                   2899,14232,4191,5790,11909,15153,1771,14695,8248,13340,2085,1166,12121,2804,2076,
                   8504,12802,219,12952,13984,4055,7949,12247,14388,15671,7993,8886,1451,12948,16162,
                   2891,7595,8749,15094,13937,14450,10709,10029,12244,1653,12608,9106,11352,11231,3354,
                   6205,14397,16074,2582,9722,4725,7050,1612,10487,11130,917,9715,14451,10687,1418,
                   7014,11635,2974,8011,7013,14991,9754,7501,4210,3395,13099,13693,7840,11236,7599,
                   9465,12251,9141,10476,8550,12187,9256,5795,1671,15726,8395,12795,4307,4080,3010,
                   4776,9609,15562,5690,8335,5309,9953,2637,866,1816,7360,13495,7415,7343,1213,
                   13792,7278,1530,13968,7352,4311,11767,1702,4278,387,6009,14276,14094,11177,1392,
                   2861,12449,9168,4117,8589,15000,2074,1934,2216,5982,3339,1390,1725,708,6126,
                   541,5487,10104,264,9584,7871,9053,3709,5760,4207,4067,3133,5577,11052,1191,
                   9877,9474,13256,9080,7282,10371,5886,12175,12973,2487,8866,15716,1231,13684,12777,
                   4778,7246,6407,9334,15911,15612,13821,4918,6055,14955,4177,9769,2773,9349,3628,
                   6412,2218,8212,13330,8393,3856,15693,6321,15707,267,2873,16259,7691,9100,5588,
                   2785,5384,8813,13776,2241,12866,3180,5112,15159,15390,13543,2011,14316,10322,7891,
                   16372,704,12962,10526,395,12359,3003,16309,14563,13674,2777,12078,6719,772,1208,
                   9230,15103,724,8552,5850,733,4815,8460,8790,1731,11765,8481,345,8298,10412,
                   7311,11858,13653,5295,13625,1865,6442,13717,1370,14857,4506,3787,13023,10947,6688,
                   651,11214,9574,7320,5558,7519,5475,13170,14321,6579,13124,2028,4539,10057,3085,
                   13698,8459,11952,14432,14467,7359,10644,15140,1968,7581,11087,8854,3336,13562,3964,
                   10632,1886,2376,13496,5638,15358,14218,13757,9757,12928,6689,10904,15256,12182,5456,
                   11168,8585,2847,12552,13118,10085,15194,10153,12140,3546,2878,988,98,16292,9632,
                   11921,16363,9363,14329,12208,10360,270,15251,14128,12253,304,12542,10066,947,11705,
                   10625,13112,4509,8003,9311,10504,2025,12371,161,16027,4493,8361,593,5036,15719,
                   11292,7222,9515,15124,9990,6074,8207,13239,4367,1593,4140,2942,12304,3689,11249,
                   12594,8142,4901,187,9041,9427,9727,7213,16131,14847,8078,8565,11730,8416,16140,
                   16281,8592,6597,8062,8387,14810,2923,12288,4598,6105,16037,11954,800,8492,12901,
                   6187,8566,9284,7813,15014,11664,4968,11408,1251,13428,1786,10799,5576,2946,5621,
                   6345,13898,2285,14359,3514,7898,14667,7886,7115,2755,11439,852,8586,5875,9619,
                   9307,12487,7969,12619,9176,12285,6638,4423,1932,12119,8400,9024,8452,12550,1661,
                   7580,10931,2337,6734,11813,6199,2707,6878,11277,5471,8628,7397,2676,11528,12655,
                   3664,7118,12214,7242,8270,13262,3971,7053,12013,6850,2571,13460,11940,15927,8337,
                   5455,3726,3759,2766,5203,2095,11581,5326,14494,6022,13065,14714,8950,4942,10705,
                   10486,3647,16121,6543,6909,13939,15473,523,8269,10422,13000,429,15376,9028,12349,
                   16357,3376,69,12077,3361,3877,14263,11243,5399,8135,13127,8033,14008,12181,13225,
                   13832,11660,5429,13933,7438,18,1183,10951,5457,11485,3289,2049,13970,8848,12274,
                   14095,10769,13287,12857,3783,7125,3850,15711,5298,14157,8225,4681,14473,7488,5169,
                   9301,13291,10179,12219,402,11716,5228,13449,3296,13182,12560,2589,11857,162,13451,
                   2542,11456,5658,3004,775,14118,14614,4986,10907,650,2666,877,793,6626,12598,
                   10308,3828,2190,8085,3701,16095,4698,2910,6362,3355,10694,9062,15287,13633,9431,
                   10724,7598,7407,9924,10208,9653,14262,11153,7860,16082,7200,16001,12595,11010,6697,
                   3979,8569,8974,7706,16015,5985,1309,2357,13744,11805,9269,1016,8640,10255,11585,
                   568,7374,1245,11623,9558,13455,11549,9128,14481,12027,5470,11094,16350,480,1902,
                   11628,7902,10306,5805,10317,12161,15660,689,12821,3981,7387,10996,7223,8829,4686,
                   4286,363,8465,5762,9136,1560,4043,7401,13515,6794,14552,9237,7865,8190,2365,
                   8745,3478,14659,13762,10295,5604,1551,10239,4695,13687,6692,7289,12979,11869,11902,
                   7614,1359,674,3634,10195,2576,5193,8711,1138,13218,2063,11787,5218,145,7285,
                   6192,2227,3861,5162,9900,9483,4849,3369,7181,5007,9434,10693,9107,4161,9253,
                   1533,9513,14975,2511,8365,2214,14577,6488,10166,4196,4437,5417,13491,12173,2170,
                   15200,1235,3725,2392,7937,2043,13916,13856,16255,5372,10619,4167,6804,2146,1042,
                   2333,5330,14723,8620,4383,9562,2250,13651,4330,1929,4015,8145,13279,6143,9234,
                   13280,5157,9329,1694,8768,4477,5991,11048,1250,12897,12177,9829,8596,7708,9501,
                   16250,7132,13282,5227,11894,571,6330,13982,8601,1759,506,8723,15714,421,10395,
                   13992,3925,8540,7522,5525,14405,7186,853,11066,12909,3919,9955,3459,7060,3763,
                   2440,7560,6586,2476,7776,6875,10157,9881,10040,14767,11207,2543,13858,14743,7318,
                   1084,4354,10385,8772,9835,12093,3230,1306,9843,4546,12590,14419,4242,12671,14399,
                   11481,2079,11796,12156,2078,11476,7530,12562,3288,11170,8818,663,8803,9207,2052,
                   8643,14759,4882,15402,10461,15268,4782,9443,3073,15545,15057,11831,4391,4842,10089,
                   503,1909,5943,3054,6025,9138,14725,7687,8771,493,4710,15852,2716,12816,5397,
                   760,2103,8608,13360,727,4232,2557,11099,2677,12265,10155,13038,10318,15622,6359,
                   16294,13748,256,12122,6000,7027,1398,1747,2179,667,7404,4716,9129,11272,9416,
                   245,7784,12185,7601,7316,4341,5684,8474,6086,7896,15209,1145,15134,14687,5376,
                   12,3707,2973,9861,3773,14204,9345,6018,8469,6835,15004,4046,1483,5282,5327,
                   11122,5954,5853,10254,11265,15180,9157,12341,2731,14039,16030,4251,6568,3433,5217,
                   7030,12947,5317,4402,8138,5599,3848,9297,7618,14275,4504,8816,5158,7768,5642,
                   6976,7820,13346,8284,12426,15550,12760,13808,4619,1573,3291,1244,11269,14517,13683,
                   14380,5556,11281,1903,13838,3615,3612,11963,2975,10712,12745,7366,15404,9859,2807,
                   14870,12090,14821,5926,7195,4109,584,4499,9871,15407,12846,6135,6239,15770,627,
                   15331,2868,9392,4958,11162,5428,955,1005,11046,4969,13526,12206,3995,10034,3375,
                   8811,6557,4494,9989,13143,12471,12911,13192,4684,1859,7325,2492,5080,13796,13521,
                   9225,5923,16177,889,9356,3287,2758,13904,13271,9352,13204,4801,3838,15833,5440,
                   9631,366,5467,10624,10980,13502,4774,16376,5931,11879,11752,9992,15467,4965,3577,
                   11196,5229,9800,2318,15558,7497,9152,9693,2568,2000,8103,1663,15701,2859,11023,
                   8564,13810,5652,14526,12132,13306,6034,16213,12998,358,2129,15728,2631,11847,13555,
                   14627,14547,13028,4562,14271,3316,11711,11878,1604,5107,9605,13814,4622,5833,12596,
                   4308,8159,1260,8480,10886,1703,10762,7087,536,9240,3673,14138,14565,5185,15078,
                   9217,9056,4266,15866,9879,10253,15869,14608,10474,7444,2062,11337,1405,2621,8009,
                   2394,14531,2906,12600,6669,11478,12157,3335,9776,8992,12894,14567,13212,9268,11260,
                   8962,15592,3833,12501,519,9413,6198,11090,701,1269,2617,2993,11937,11932,3240,
                   30,2126,12272,12008,14182,3238,2647,4609,640,4390,11502,9720,14568,4837,13297,
                   9403,10580,3496,6099,1293,6615,6885,205,4612,4643,13554,11744,70,13662,7773,
                   12770,5822,8219,3597,14508,2588,11203,10892,13652,15837,2229,13567,8082,13974,12714,
                   3237,1340,11903,11324,4218,2990,9654,1948,5058,6590,9601,15338,11753,11710,881,
                   1588,15290,14395,10198,9354,5754,12051,2465,899,16045,2018,2892,6787,11420,570,
                   14663,4335,14660,9583,10621,15476,11325,11868,13244,10531,14728,3900,5791,10655,2926,
                   13092,1761,8506,7758,2117,3690,13731,4404,6749,16362,10966,12451,1860,15659,1388,
                   15144,5435,1797,1233,15542,6978,11819,11936,416,230,11933,11818,4295,8233,11113,
                   13461,2734,7258,671,6388,16010,5407,14579,5660,5305,12083,10923,8458,11037,16036,
                   3728,16113,12514,8090,6791,5361,3613,11633,5390,2781,1669,4392,654,5617,5628,
                   4715,14523,121,3261,1884,6860,14746,6337,2997,2238,15657,13414,194,1584,15137,
                   9486,13869,6818,777,7099,12871,1061,15086,12380,6030,1290,6100,3697,16358,5770,
                   2797,3513,13840,3859,13409,4799,9796,11824,14183,5060,13576,7052,11109,9130,8051,
                   14787,2474,5383,8557,5270,8500,3558,4862,4357,332,14480,11275,4954,8706,10118,
                   13573,278,10553,7642,652,13499,13671,4672,9492,2685,2987,1960,13976,14235,14006,
                   15982,6493,13304,3123,5755,11887,16078,9187,2809,1311,8040,5016,6886,596,13644,
                   12702,14863,8798,15595,1178,2619,14300,13517,8654,15324,6245,3840,15858,6902,13481,
                   68,11149,10872,6718,4346,4551,5304,11951,446,5031,2314,3228,13246,14206,11642,
                   14820,3231,11466,4273,8325,5140,8738,7534,3855,2162,1542,6434,14197,1581,14764,
                   1020,10488,7477,4077,5412,8355,2145,14414,1194,6343,9849,7390,8401,11080,1167,
                   10663,11539,257,16178,16342,14931,4797,6313,14927,6451,12373,11735,14527,10159,4560,
                   3731,5449,14985,8332,10959,10152,13854,12863,1552,15072,8953,2994,14173,9004,12706,
                   8054,7725,170,1840,8542,11479,11797,454,12309,15661,11286,3061,5378,12774,9746,
                   15098,12189,13265,6760,3152,5842,13490,11369,12972,10808,12896,11411,2838,6133,14009,
                   11159,10949,15257,7785,11553,8551,10731,15099,12167,7143,3370,3826,2309,15678,5809,
                   9461,10539,13630,5866,13647,15246,8356,12941,14915,4802,11667,13527,10970,10361,14252,
                   9282,3097,7384,11103,7119,14348,5411,403,11194,10220,15621,9411,4034,215,15456,
                   10495,8830,4659,5147,6957,5657,15327,2948,6252,4889,10030,5062,13268,15029,5200,
                   13135,7039,51,10689,10028,7948,10673,15723,15689,9464,10727,14129,10975,9027,13220,
                   1189,4406,8390,14097,3226,15673,6732,4747,10154,11530,13800,7524,3119,14653,5826,
                   16246,11823,2127,11175,8849,1262,1134,8115,1385,12354,6148,9789,3954,6639,11076,
                   13410,16291,11033,2922,16132,1709,6698,222,12431,9738,13789,7909,14848,4909,4669,
                   3031,4497,6258,11008,3688,10485,14515,455,12159,9260,6954,12782,7509,12812,124,
                   517,3732,13214,12445,217,6211,12765,13227,3331,7951,12735,12467,9089,14712,2983,
                   7189,520,7344,14489,7824,7280,15146,8742,7413,2730,11588,810,13910,2438,1728,
                   3068,5049,9029,11145,8242,6642,6975,2454,12280,6149,12773,488,3002,10866,4691,
                   8435,4997,8130,10012,2670,8456,16266,7575,5450,160,10988,6450,12131,14257,3274,
                   7832,8599,10522,6923,11994,6031,9832,13070,13319,7723,3642,4313,3053,9199,2430,
                   6572,4595,3711,16333,15790,5906,1403,14216,13469,6948,4640,2645,730,6570,2634,
                   6206,1749,7198,9918,5348,14806,6203,13141,874,3483,1518,15788,2264,414,108,
                   8560,14897,8980,15589,16367,11615,8285,8764,15012,9739,12294,3617,1937,14642,1019,
                   2064,14085,6325,3027,9784,15740,3652,15300,13215,12319,15438,972,9169,10772,1861,
                   11922,7399,2429,10267,16234,8880,15785,14371,9346,10210,13310,8226,7533,8613,9688,
                   12734,12327,4527,7417,12910,11676,3663,3717,8311,3928,3067,5679,13539,1255,7196,
                   13108,8439,10231,8036,6102,7968,11072,16335,7122,13746,2014,14581,1803,3150,8149,
                   4660,427,14574,681,3832,11809,10516,2360,6117,13308,2444,1517,9448,13713,4689,
                   3156,15267,6283,11958,8091,14886,6063,2248,2398,4671,3891,3303,8801,4060,1993,
                   7977,8531,8665,15113,2815,6598,14778,14837,2317,945,9914,5046,3898,5009,16289,
                   2006,10977,305,15204,8462,487,9596,1472,4638,11084,1660,10954,13119,9294,14951,
                   16341,3906,9937,14259,11201,13183,11483,7531,7633,8797,14929,16183,7641,5280,10574,
                   7740,12754,6891,14411,6940,12970,7726,397,13255,9567,16370,13293,1096,10125,13766,
                   7966,15307,12639,2854,11471,4547,3982,9750,11011,11248,11760,4309,11220,10309,11794,
                   6668,6868,5245,2037,16057,10175,7095,10691,1652,4592,14812,5284,1843,12633,3618,
                   13884,9823,9177,11074,12757,8704,15514,12840,7463,6069,6064,12903,1172,173,723,
                   15176,3619,12614,8879,2602,15003,5358,2855,12588,7853,754,5419,7713,1871,2044,
                   8001,14403,1513,10279,6219,4129,13007,7481,3665,11100,13826,9772,3869,5388,5711,
                   6318,14702,10326,12891,9670,2967,5788,10094,8288,14398,11474,1498,8489,5989,13721,
                   8630,4365,12914,8538,1892,8702,13058,2198,8308,2592,13704,13534,14596,10583,5528,
                   4571,15813,7585,1153,2565,6914,1912,2936,1876,1425,530,12061,13645,15988,15585,
                   12150,8055,3341,15511,8752,2255,110,9288,11865,13975,15522,6968,13478,5342,2713,
                   307,6422,8004,14287,6094,10126,6083,7988,2386,3627,1331,1682,14111,12466,12326,
                   4913,15591,7136,15239,459,4006,647,13229,7367,11636,3413,10507,13966,12860,2723,
                   1381,9149,3883,12572,6890,8705,12620,15430,15947,11617,15551,9669,7182,13226,12322,
                   7215,15861,8783,13399,11851,7772,489,12356,12164,9747,13685,10815,335,10519,10359,
                   4446,12312,7508,16287,2451,2831,6424,7765,4575,6799,7483,11,13877,8394,10737,
                   9037,5289,9791,8674,10264,13641,10667,8505,8903,13026,14486,4933,1825,8697,15163,
                   5464,12314,125,5409,9557,11519,2717,15892,5963,688,11289,14827,14905,14086,3400,
                   9527,5186,628,8833,8330,3092,13964,5328,1597,885,1999,603,4535,15587,12623,
                   15515,5207,4438,6361,5427,11651,15406,15064,4903,1415,10482,3651,6405,7980,10381,
                   13286,11179,6876,12913,12749,13967,13855,12143,4719,3135,10851,2240,6051,4325,7098,
                   11991,15817,6895,4009,2405,781,7176,14838,3268,13197,14937,15501,4332,14185,2741,
                   932,3248,9425,15964,9671,12664,6530,2884,11801,8993,12176,11410,13837,6717,6186,
                   11040,6065,12627,3065,4757,14445,14170,3918,11440,12470,11677,6877,12859,12678,8539,
                   4946,4515,10082,7299,6690,2172,1098,10068,3023,572,12944,13492,10945,9756,7000,
                   13332,3353,15433,3311,10601,9629,12966,975,6272,8357,12203,3682,7848,12926,13493,
                   7031,11597,10679,1450,5303,6565,10669,218,3273,4703,8372,5035,8442,3264,2955,
                   10469,10863,705,4375,15189,12937,9628,6962,7175,12576,7727,12174,10809,9650,4956,
                   13328,4429,7288,11323,4656,10049,8635,1602,15638,3196,13734,10542,3520,8261,1101,
                   9074,7557,2034,10388,3953,13272,10276,11739,16212,11141,10423,465,9002,2101,9635,
                   7480,12652,2111,361,347,14986,3308,3713,7770,6518,1772,4578,5214,5793,4624,
                   8273,3786,10903,3661,4472,12805,8902,11748,4563,13040,4205,3962,15219,9457,2187,
                   15178,7427,11532,10319,13030,4204,2984,9507,10640,5042,6810,14151,15597,1253,8728,
                   14792,8495,3578,104,14664,7607,3390,12682,2199,6446,6256,10115,3141,14715,11126,
                   3460,5748,15610,16248,12383,9833,7555,9621,15913,1675,8045,14762,4820,4227,1324,
                   9010,2449,338,3454,2206,5567,7295,9910,10219,7369,13849,11911,2927,2956,3142,
                   7429,9015,3394,10721,3564,14289,1265,13202,10282,4,14824,2495,12481,7197,1763,
                   5941,10982,4508,5836,2632,3624,983,10955,12553,424,2371,8267,3315,10916,2029,
                   8032,11156,2651,13241,15210,2901,15756,15040,5201,12241,13445,10435,2125,357,6202,
                   12413,9988,11675,14866,924,9886,9480,6778,6823,8536,13813,2871,8313,83,328,
                   7160,14159,14192,8870,393,7077,6674,1921,14440,2980,3620,4738,4972,13802,10913,
                   5474,5724,15553,9975,16043,9812,16147,15984,636,13584,3897,11200,12561,7167,1609,
                   13901,9275,3362,5828,8834,10171,11678,4685,5514,1476,14936,12880,1407,4115,9135,
                   3139,13103,1264,11696,4800,7998,13587,2200,7900,471,3977,11803,14566,12318,12444,
                   15761,9205,11335,1139,12255,9026,1715,13893,13833,11160,12764,12323,646,12743,13569,
                   411,3253,8445,15483,13959,928,14649,8206,11003,2650,13129,8721,1979,11904,10530,
                   12088,14207,934,4091,15865,7877,14280,1755,396,12579,10803,9475,16058,14956,7616,
                   9943,11106,3970,6761,12168,13299,1524,12238,15028,9353,11694,12996,10277,7553,8961,
                   14211,3865,6142,11398,11401,9235,11418,5226,14910,4944,12856,11178,7409,948,10178,
                   11192,1097,12582,3095,15906,4836,11835,1525,13266,16100,7803,9059,10190,12048,3122,
                   11736,6035,12505,6116,12461,10211,5152,7268,8967,77,290,6229,7722,12384,9698,
                   2331,3575,14362,3081,869,5022,3601,12976,4428,10834,8392,12931,7001,15874,7450,
                   15037,10491,13608,5813,10660,2084,3831,1819,14748,7873,11613,7821,6581,787,960,
                   4847,5319,7835,15899,5337,14774,8297,9372,14446,11524,726,14802,3120,3177,13588,
                   17,16380,5165,14021,9390,3102,8485,13384,2718,6335,14189,5086,5473,2168,6460,
                   2197,9759,2213,13373,8484,6843,4158,9831,7659,1326,4871,1989,941,5625,9764,
                   6146,9564,8782,12769,3818,2705,807,6108,986,15374,8291,16283,3858,12005,12286,
                   16290,3233,9091,11982,195,7009,2500,3705,1899,10454,14264,10623,1142,101,3518,
                   10515,842,11050,1787,4663,14372,6918,7838,15120,7526,13750,4952,14109,2417,969,
                   7233,14719,5462,10434,13136,8804,8549,3297,11198,163,11205,13952,15536,9559,11271,
                   9238,10227,7241,6582,11112,11941,7230,3806,6131,6453,2373,14732,14217,12399,1168,
                   14390,1795,1520,5114,1454,2837,5354,12718,5343,6903,12075,3494,14054,9432,1334,
                   490,7251,14632,7025,12172,11368,12927,12945,7414,10752,10939,2377,13670,12036,10564,
                   8092,11706,4775,7154,15509,4636,10458,4089,14994,3326,4000,1707,5718,6795,11304,
                   8655,12068,5262,4258,13797,11685,6632,9124,10214,6287,11666,12207,2520,8616,4183,
                   4431,7346,1072,12687,13705,8223,2397,1254,12478,9916,5736,2010,10856,6943,9938,
                   149,2599,8941,8988,9368,8349,10160,14650,11846,11745,6574,1778,3411,10467,16369,
                   9602,10934,3965,9548,4491,8083,11862,410,13230,8067,9286,10119,12031,13595,1141,
                   12011,5061,16164,4458,2680,10007,5980,7227,13180,3896,7999,13207,13365,3176,6757,
                   3415,4036,1798,1140,13574,3741,8670,6395,15531,16311,643,13923,5209,7377,14888,
                   4788,5242,13338,5812,2083,6841,9083,8447,15763,5051,3529,9705,2538,4839,6523,
                   5986,7075,60,5294,10895,7583,1280,9121,13715,12198,5867,9430,11234,3768,242,
                   5994,14199,388,15889,10265,12801,8397,1554,12060,12703,15247,12200,10339,5594,2251,
                   11393,11859,10893,16102,4745,1689,4948,9724,1579,7253,664,11849,71,7800,5637,
                   8715,6013,4234,1591,13498,12037,3720,4591,10870,2776,13956,2466,460,6403,1041,
                   6167,14516,11625,10814,12776,6693,11320,14603,1623,16180,14753,7841,10722,8784,5562,
                   7710,7,10921,3084,5555,14107,1285,8154,12686,13535,4819,14780,514,5901,9594,
                   15343,9449,12509,9120,13629,1371,10898,8253,2835,5988,12675,16108,539,1791,340,
                   9321,6249,1304,5681,3691,11917,10611,5974,12986,10543,6301,6246,2622,901,1192,
                   10032,255,10111,11259,2356,12490,2015,11537,16295,13436,4953,6429,9102,6456,10062,
                   14219,10943,1353,7639,191,15491,11314,10294,9778,5896,12585,10124,102,8925,5921,
                   2587,6029,16081,8971,4605,10849,8812,9494,15921,15048,7767,15023,13881,353,4254,
                   2770,2268,7908,12296,15109,4811,10756,7279,7033,2151,11684,13520,4147,7313,12266,
                   7525,13169,4973,6037,7681,6740,6989,11618,4618,11732,5653,8537,13151,11757,9604,
                   3271,5297,14238,14768,4919,10822,8068,15945,15806,1176,12656,9773,6348,5873,8605,
                   7273,11161,13224,13981,7336,6716,12898,11630,3614,12003,3512,7002,6744,13996,1122,
                   14860,1900,7368,13091,10139,2865,384,6945,12142,12862,11378,16254,11458,14742,5054,
                   509,7235,6217,15497,15786,16274,1628,9487,11987,2089,2066,4532,15355,9873,9201,
                   10,12793,8064,14425,15022,13783,7205,1559,12616,9822,6772,299,8929,4184,14639,
                   8254,1714,13223,10391,4100,6200,5291,11057,6344,9274,13186,3563,7565,11693,2759,
                   1846,8449,14890,6844,12343,811,2828,5074,6115,9319,11377,2042,7111,15527,4143,
                   7934,5208,13602,6484,9730,3587,8237,4554,7629,10447,7904,7439,11164,4468,5606,
                   15095,10685,15472,11136,15494,4328,2555,14620,2574,1277,8657,14618,9962,587,6176,
                   7090,13452,15537,10532,16186,13676,2467,15482,13235,3852,5038,10081,3383,12832,5329,
                   12748,12861,10759,1531,11173,2048,9160,8525,11864,12715,12043,1961,14550,15363,7337,
                   13834,11423,6331,10670,4054,1690,2690,10197,4048,16325,9748,11431,10394,10133,4722,
                   13844,1123,788,4024,6465,4544,14379,14901,6921,6532,12045,14234,11158,12180,2702,
                   14676,1939,6721,3243,10378,9923,7147,6708,7411,5164,13369,3224,9450,4005,4791,
                   14028,5949,14026,5948,8420,2167,15680,8725,7157,15198,7029,5531,16031,11590,8160,
                   10165,15831,9552,2433,1373,14720,1732,16053,4489,14457,7314,10649,3774,13483,3495,
                   2765,10086,7018,14716,5798,10635,6473,8382,1075,3542,6897,4170,8263,4152,8110,
                   8563,15917,7149,8555,303,25,5782,6121,10401,3247,14492,9836,15803,2065,12437,
                   12824,3401,1489,1131,16117,16089,15382,5746,10768,11176,8391,12259,15487,10224,5351,
                   4022,8455,15275,6006,790,5554,13701,2416,13438,1683,12733,2426,14830,10595,14556,
                   3404,8622,11211,774,5722,4881,1881,995,4432,4148,3450,6678,10974,12252,15742,
                   528,8414,7418,4635,6266,9171,2409,11772,14564,263,8473,10129,2462,4467,8515,
                   4867,7023,8767,5694,6811,13047,196,5756,15253,3843,5299,11185,7161,13157,1894,
                   9663,9018,5953,4050,3325,8986,322,16013,1186,12907,14444,9005,12148,5884,3186,
                   1627,1466,1537,3462,14622,1175,11825,12009,2740,12884,8701,9012,5087,13376,15038,
                   14640,13158,8871,2769,4056,6435,12103,5995,13637,4829,3936,7928,6672,11571,3772,
                   12089,13247,1011,15938,3864,13276,1611,1507,4389,3322,12398,13468,10942,13756,7763,
                   14794,6959,7328,7942,1247,5142,6553,1377,6411,5532,7452,10652,4190,14007,12044,
                   5551,9884,13818,14769,9767,7378,737,9802,14917,4029,8167,16156,1891,14939,14327,
                   16124,12210,9283,1563,6439,3275,12374,9936,12559,3572,2502,11242,11152,13421,10455,
                   15772,15796,1704,5510,3317,11750,6369,9827,7619,11605,10767,6008,1300,9972,13252,
                   1754,4380,5323,9396,7402,6095,12724,3565,13101,2507,15196,4961,3881,14657,14823,
                   7958,4679,14685,607,12067,2618,1987,3113,1241,15521,15459,8659,6752,9273,7754,
                   6681,16270,5013,7017,16066,10858,10323,2366,14876,6578,10914,7079,10599,8241,4193,
                   16125,14250,9362,10969,3305,14976,804,3013,6592,10456,4336,10172,4426,4394,8316,
                   1547,9742,15318,2059,1882,10113,3835,12216,5410,15221,15455,15111,6537,390,837,
                   3798,5000,2284,11059,1684,7036,13323,3574,15052,15676,4834,9904,154,14536,9347,
                   12458,13431,4662,7202,1738,1491,8856,14900,14002,11626,5557,3638,4168,15642,15746,
                   9694,1574,10674,15670,13471,1169,6240,1452,15291,11883,6204,10697,12670,11475,5623,
                   15721,8000,12647,7187,11436,8516,6667,779,7945,6941,12574,8862,1811,12113,2144,
                   9535,4794,4243,11472,5198,2535,1401,635,8065,13879,5509,3556,7930,3911,6383,
                   8982,10924,14466,1673,8931,5065,4927,7245,15651,13164,2981,7612,6409,14171,12906,
                   13359,9373,2908,3040,10686,10708,10639,6677,14502,2668,7315,14050,4163,8545,6731,
                   4754,9550,16184,484,4999,14433,10925,3108,8257,6931,10109,7489,11188,9490,4441,
                   3158,9896,142,1328,12026,11274,6729,3182,5552,9182,12806,4932,7825,12334,7219,
                   10131,14081,3246,11124,6023,3279,8991,2282,6589,8916,10122,14454,2669,9069,7792,
                   6830,6352,11855,3596,15637,2047,10418,1286,10484,12307,13682,11624,10102,1469,9678,
                   3985,120,11972,2560,4445,11734,12133,5167,15685,2907,11792,5174,505,9210,14817,
                   14369,155,10289,15534,4536,8508,9622,9299,4302,14558,14626,11747,9946,15050,13978,
                   15362,11306,9236,3915,8957,14115,10594,14545,4303,6168,14,16308,10869,14139,11773,
                   13213,11802,11833,9721,5670,4455,1078,10053,12498,680,6489,11362,5661,11948,1802,
                   12492,2749,2595,4030,4712,9906,15117,2783,863,15278,4413,1087,8368,8200,8973,
                   12688,10582,15130,9031,1601,5518,1622,13688,3213,10148,15629,4084,11783,15868,1049,
                   2119,15808,15258,11212,4987,4931,5945,13947,8656,13943,2554,14180,1174,2073,2352,
                   14546,11746,14672,8979,7228,8327,13488,7024,3800,2244,5730,8709,8255,13890,14191,
                   15039,12434,1018,3256,16151,4132,6629,929,13237,13553,10161,3118,12269,598,2303,
                   14822,14294,3479,11313,11898,9582,4334,11896,13055,105,7887,11062,3811,2857,3464,
                   2746,14628,8978,6990,7548,14011,2703,1343,5973,8340,7084,1701,8304,606,14298,
                   5377,11564,14903,15649,8997,4934,6766,10076,8249,10658,4096,3062,10005,1753,15429,
                   3922,12662,10327,5380,8108,2155,8096,9444,5495,8048,2246,12329,9088,11127,13064,
                   14059,7019,5463,13442,14046,1733,8621,11388,7686,11512,8841,4897,11906,3901,644,
                   6650,13467,2372,6372,6827,6924,2932,6545,2350,555,8427,13859,11459,8112,269,
                   11977,6861,13344,7872,9021,7544,16181,13691,6802,9577,14833,2262,4883,11492,2979,
                   7045,13077,8044,12105,1580,10041,11455,13819,14239,1548,1823,1990,9762,13356,8296,
                   1056,7163,12532,14836,13707,4818,4924,1649,7913,2181,2475,12016,10646,3508,10027,
                   14804,13051,8729,14221,7762,1214,9358,6226,5236,2021,15617,13362,3121,14791,10026,
                   12411,5349,5773,4359,11031,8386,12611,4593,5619,6026,9211,14535,6644,3014,12091,
                   11643,14656,14295,13106,2494,14904,12822,6747,8380,14113,2427,2263,14756,14971,8058,
                   14779,12533,12878,3269,9821,9455,4963,5004,16171,5613,8079,11020,12298,4908,4263,
                   976,16260,1445,15191,5340,4507,10900,6548,6789,13846,1901,8799,12062,8626,15446,
                   13144,925,16159,7422,11641,2806,1460,9280,3498,5268,14319,2367,6966,8937,3418,
                   5844,2135,444,9818,15818,12516,6062,13605,7376,13908,6845,248,15018,9593,7464,
                   8981,12422,9509,15902,14378,14003,15648,14688,14826,12823,10479,7883,10098,3456,13284,
                   4945,2989,8747,4803,12204,4028,14244,16298,3606,1362,854,4720,6145,3034,9147,
                   6312,12129,16182,12566,4796,12126,129,7782,1765,3986,13196,12881,1890,14249,10018,
                   10092,610,4012,828,16155,619,1699,1273,15261,9295,12555,2038,3874,6054,10825,
                   13259,16059,1944,9341,6503,4203,14999,4858,3399,16145,15066,9151,9229,4083,8059,
                   14834,7856,7434,2510,11358,14331,3304,7236,3686,4807,2301,8211,67,8333,12138,
                   13011,346,5204,9935,9755,10716,15426,1508,13509,4088,8258,5133,4859,14962,10776,
                   2075,5359,12636,11576,4047,7655,1155,3771,1631,3320,9276,12429,8765,11045,7812,
                   15062,8893,14893,249,15480,10560,13880,13782,9165,15452,2192,15271,13269,12239,9094,
                   5708,5027,2159,5321,8618,10490,13336,14190,14641,13133,15757,8985,8012,5717,7851,
                   2762,8251,13780,7766,14549,9947,14364,15677,16297,9223,15544,11501,2149,9419,5741,
                   4157,15016,8892,12848,4902,14966,9150,6049,10281,1927,10578,12145,1553,1783,8730,
                   4396,1983,11775,5184,9142,5869,5130,15170,3752,3824,11993,1060,16110,15745,4510,
                   15725,10605,3283,10684,13936,16008,614,12166,12188,2662,4772,9231,10877,4480,6270,
                   6637,8650,4810,13790,6536,14352,8664,12529,6496,5482,9907,14587,513,5768,13434,
                   7527,9957,4611,10999,9514,8057,7459,1781,8245,14598,9030,2795,4344,11563,1144,
                   1585,11985,9866,8583,10928,1969,3817,250,11926,5434,12337,7281,10372,6800,6184,
                   321,1770,10656,15749,1206,8876,15733,15391,10854,5543,9806,5465,12810,8353,4885,
                   6813,10589,7906,4068,15083,5131,535,5421,9883,3845,12631,722,13036,7426,11586,
                   9156,4461,1249,463,8944,8410,9126,4374,12965,5341,14854,3589,8408,10957,10084,
                   14291,2506,14035,7156,11371,2171,5777,15569,12544,8463,15696,6933,7897,11561,13130,
                   2900,9406,436,6528,10070,1410,5513,3963,13033,15454,14350,9912,4145,7221,8858,
                   3204,2753,5663,6392,679,1225,6630,4742,4971,4058,5802,9009,7137,12739,714,
                   5573,8053,9401,3667,1848,12201,13646,656,1201,271,10973,3842,14154,9476,5960,
                   10948,12183,14613,15809,1272,14949,9825,7794,4398,6780,6282,12512,11496,4783,2193,
                   15027,3350,3945,8454,14103,676,551,14590,4412,10353,2965,6284,5854,6017,557,
                   9063,11233,4990,8,11882,14394,5264,9016,9809,1966,15754,8182,9733,3510,12443,
                   3653,7940,2541,3048,6995,7967,12587,577,5129,7503,7730,10452,3173,4887,9888,
                   4915,1896,14343,9743,9191,6197,3039,15606,12070,6244,2949,12232,3125,3218,2869,
                   11656,2952,9370,8230,8419,2528,6278,11877,9600,7954,15800,9595,13711,2278,937,
                   10441,711,9221,4979,822,10189,10573,1465,4533,13873,3958,8913,10941,5639,3018,
                   273,14551,13979,7788,8521,1946,15572,3813,2625,1829,1162,7362,336,13405,987,
                   11143,428,1421,5221,8129,5230,14092,5747,448,4929,10192,5819,8999,5825,10855,
                   15158,10613,546,15851,1745,2324,5250,1974,672,10442,856,11494,10460,11638,9858,
                   12847,11650,3490,1092,1344,10500,5627,1712,8007,2375,5707,2184,4750,3424,6848,
                   4368,3,8736,2709,8873,14992,1509,3923,14700,12758,15946,3352,12933,3551,3894,
                   3001,7786,12446,973,8205,9985,10177,9555,6659,581,14865,8627,8820,168,6076,
                   3681,15025,9164,15220,14351,12225,214,8658,14306,16326,10259,3751,8423,4920,2615,
                   9993,11713,8209,10520,4194,7046,13938,11137,10493,224,11901,10620,5155,5096,15020,
                   10561,13958,13234,282,7579,10225,14098,452,107,190,13761,2483,7153,13940,4329,
                   15787,13864,2152,8163,4333,12882,4893,9586,840,10042,4517,2460,7155,13505,3340,
                   12709,9462,5260,12622,12841,5957,3523,1058,2097,1240,14305,12716,6969,16068,112,
                   7110,13919,2287,5310,6394,13599,16197,2548,14539,10288,13453,13953,10290,7510,6507,
                   6617,11930,6979,15056,11500,5925,141,1484,7049,11616,12761,5725,13173,3437,10091,
                   2293,8403,11720,7496,9902,7350,10743,9608,16139,7973,64,6379,5776,15203,6092,
                   1676,15367,1947,1500,9422,7682,3893,4260,10237,8534,9159,9084,6223,15989,12705,
                   4534,12839,16366,12424,4912,12737,11807,8963,1179,12064,1252,13048,1851,16169,6832,
                   84,2818,4410,15699,9489,15323,3038,495,4582,13068,16249,10821,15910,2354,7610,
                   2020,14801,3190,620,10221,12221,11534,6358,16242,56,5522,8034,4085,14606,3452,
                   3555,2434,2655,4646,9814,2046,14510,12984,3197,5806,1274,14384,15747,15654,5144,
                   311,15940,14902,14689,7244,14439,10140,3755,15644,5145,2239,11981,1389,11924,11287,
                   12160,3595,5965,6188,5750,4299,7528,2659,8807,14389,10675,3227,12261,4759,742,
                   14365,15053,12194,5808,14032,8724,6846,226,5166,14529,903,95,15722,12249,2678,
                   9976,3857,10837,5111,6970,15206,6932,9488,15604,2858,11728,16195,1076,9048,6441,
                   6320,10839,4110,4793,3851,11183,7486,5021,11428,420,10812,1230,5037,10995,5622,
                   14401,15688,12248,4511,15091,10735,1670,11742,2630,5654,4731,8877,15157,10216,6311,
                   1226,9408,146,10627,12441,9785,14130,529,16111,15089,14385,15643,1207,15154,10274,
                   2267,7932,6212,15296,8183,13132,15041,3795,2456,9204,13216,5050,13614,5239,6032,
                   16188,8300,114,6524,11654,626,14266,15797,7333,8636,4693,42,1642,3416,15835,
                   2205,5430,1409,8881,12457,13865,15496,12417,1519,12395,16332,5780,2291,7604,8918,
                   14267,15773,9468,6534,15341,7955,9837,14083,5641,3805,13824,1177,14612,15259,5223,
                   10511,7584,12692,9683,9367,6894,12872,14885,9819,2447,3748,962,5860,1090,3675,
                   7392,4951,4589,4804,9553,14042,3839,11699,2204,15780,2228,11860,1126,32,4343,
                   16272,1942,2888,1617,838,10024,3046,3258,8684,1744,15394,11517,4711,10147,750,
                   7101,9659,12073,3841,7214,12767,1955,2130,7876,13250,11779,4267,14609,11782,2071,
                   4542,9869,16017,13334,7451,9855,15890,4288,3622,7651,9588,1270,5070,7112,10285,
                   623,7822,389,13639,15877,9854,12818,5962,3449,8343,6123,6080,5336,13354,1665,
                   10631,14899,9508,8788,2875,13295,3094,7670,3764,15613,10820,1674,13074,4645,10000,
                   7148,14072,2339,15931,9495,13779,3476,9324,10535,371,8336,11114,3148,16199,2338,
                   15919,6293,2904,7653,6097,6243,16073,14209,1010,15647,310,3301,1595,8069,13823,
                   15431,12759,441,3179,8606,5767,4265,28,6263,8121,8910,4017,1360,2761,6427,
                   7303,5190,9691,12889,9424,8826,1726,4377,9998,2745,1217,8882,4907,2656,2323,
                   6364,7255,9864,1023,2917,9247,12046,6492,13178,637,5338,2903,12704,15584,4094,
                   7192,9317,2572,2938,7827,6603,7970,6793,8890,7201,11247,6323,3743,4655,210,
                   5492,5714,15096,615,11946,5406,1187,14168,7707,11255,9868,15873,5895,2811,3506,
                   6124,5357,7844,16192,16216,4492,10990,8787,835,11591,14038,601,1315,717,5871,
                   11955,11036,8168,2827,4238,16315,9974,13175,2019,11890,2348,5108,8071,4704,1357,
                   613,4488,14048,10439,73,2036,12605,13258,14957,2849,9001,4606,7065,6563,4362,
                   14315,7016,15524,113,10472,3423,6242,15937,10698,2583,1479,8718,12052,9186,6028,
                   13773,11245,7861,8303,4988,4854,1339,16116,14091,6538,9641,10008,3485,4699,11226,
                   7355,3466,9794,7603,13300,7802,13654,4744,4700,5864,7621,1429,13722,538,15088,
                   15744,3729,11957,7563,4524,16088,14090,7485,3160,3646,11133,1171,2055,14251,14326,
                   3298,9636,6939,21,7212,11019,12290,1708,6785,821,6911,9839,7972,15564,11025,
                   8417,8024,2715,3398,14965,9813,13177,4305,7748,3257,14645,9716,8406,829,14945,
                   14247,8166,7423,14868,1952,9816,10680,2890,13578,4459,6783,3802,1850,15599,5612,
                   14844,10536,3267,401,4734,888,11688,12124,16343,13690,14752,14928,12567,14463,9551,
                   13955,10533,15766,8301,9890,6912,16024,16217,1077,15702,2549,15532,3149,15929,3541,
                   7577,315,8314,831,9804,5863,5137,119,3106,10368,3966,12999,11738,2120,7648,
                   16025,16193,10403,6566,7035,1228,4281,9544,7372,6608,134,4602,692,6807,6139,
                   2525,8176,3016,12455,10266,9979,4150,2310,8094,3131,3262,15624,57,498,313,
                   12271,5827,13069,15611,11416,7133,1815,4318,13857,11379,10262,8136,7690,10842,14852,
                   1444,2498,971,783,419,12367,8457,2699,1523,14312,5012,15841,4342,13866,1629,
                   5800,7697,2799,872,8593,11026,8290,13407,5506,375,2450,12784,2007,12540,13411,
                   12287,10964,9633,11536,13749,9222,15054,14918,3607,719,1065,2288,8688,1869,6625,
                   500,3938,14562,10868,642,13600,2412,5891,4239,16041,8279,2271,5881,9770,7020,
                   16364,5082,7306,9749,13990,15460,10258,2307,6346,2141,3792,15791,12394,7123,12488,
                   8019,6436,1413,3447,3907,12556,12125,16179,1422,1874,3033,9958,10273,2930,11278,
                   481,8116,9484,10181,545,3377,11146,11999,3696,4601,2402,11920,10967,16321,7021,
                   15588,12425,9603,13560,12581,9566,10861,7890,8824,1102,11708,5930,4993,1114,13367,
                   16,3932,563);

END bchp_roots;

