��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P�|5js�[`F�q�t�(���(-jp��
�����-V�N?�;�� S���H7L���S�w�Wj�K�DP2�_K�=@�%��՜��-d֥��K��8 �R��к�u̧J�'�U,��O!`k�	vR:]L?�q�`�Oم\�y�ˆ�a燺{6����/���
�C���2�M�z1S=^�J&��7�}J���b��ĥ����g�S����j�/FY��E�ݪ��f3E/��m8������RTWq�u�AmҜNh�=P�l��"������8��mi	Jm�l5�z��&I\Y	�q��H������p�hfU���� �q3�ds��okn"걱�U�fD^�z3k§/��{��^H��hQ��,�ߌ�����w�	�#߹Py<��J�$�h�m�Oq*�8��j�S;�c���D��
^}��k��7܁�6�:��^�����N.yyx�s1òQ��V߳�Ҩ���Te�]L`q��6Se[݋�x����; ]����"����)ly��hn��{w��p��t\D*��#�C<�uj���K*�gQ��p0œ�'����[��ꄦ|���F�h>u >-S��R��� ��>�+���?���	�pp��G�ȸ[7���NR��t@����h�z3ؿ�X����e���h%�4.k����N ��D:�X|��];�J&L\<zq��]��s���/�Z/ ��4>us3�PۮΟ@�������yRY�N�G��:w;QC��5��cDz��S,���BP7��R!qY���E�K3T��q�be���d��_"S_h�<KOM�,@���%��ހn7v��4�jѸK�)���.AW�6{�6�敹  �B�)�A����s�n�����.i�r�5F��V��Z�\Zm��~W�,Z
b���L�C�F5�kh�w���v��6���Ef�0A��qD�����R���*b�4�}�Ķ��6�nU]���,T��k��p�q#Px)B�;�GϽj���T#�|l[ދ|'�MbL�,Y:�EbH#��<귳�C�{��o���>O�	�e�����(�T
C;�.I�N-�!�H�֤w���`���;K����8��X�C,y.�(y"�Cj�"�t�jQ:��f��a^�_�:"�4����t��D���W�r�"U���� "���r�!�=D<�����u1�]�Ӷ�����P� �� W�7�'��F�ݴ�~�Ix��݄��Τ��2˥�[�b�?VA@(�gy紷Z���{�a��1����AM8����_c���\��Q�G١%���~$ 
�ӔH�ʹS��gG�ֱ"A�Vc�U�r�����3=zA>���D"��}�m���[�,�E�f#��yx�����x���:��结JK�\�L�G��]i�q�x�wc�d�٥W������{@��i��Gv�?�5o}�(��+�p��!"=�#� O�2ݽ4͈GS�ߵ�%�) x&1#Dt��s�dMDel��cD�6 a��U��e�<�ѻ��~}c72��4������f�g�F��A-+��:�L�"��<n�����Sɀ����;��U��NiԄ,��*4ɼ��As^�=���'cy^�a�L�y�� [i� �Zx�t�WB�~D��MQ�ޢ��άR5�b�o4�:�f�ܮ���=~5Ye�Ȉ7^D kX*q�����t�`�I��X�mX�g��"8{VMVYVC&��m-�C`��l��T�ο�J"��\L%SJ8+�7V�zL��>��U�h��c���~f?�����-[�L���Ǿ��h^��#��ި����'|�7�5=/�d�:�jY��_�5��H1����R���=C��y����c_��5g�Y�q����`�����*k�B..p%x������c�c��N��R[���y��\�YNN4~�"���Tb/�14�q5��Ir�
~�e���'��'�!�-,į�e2��^�]���%��
nQ�%y"������zI ��� J����o�U3���m�U%�n6�h�:�F�|0ӟ9#����ל0�B��CmڑZM�|�@a�Y���2�g�x��/�?ȣ����`���+�?=���5��������@me�6���l��w�ҿo~L;���z�%?�7TCT����2w�+���̗�lUp_H)����m��$���!��M���}�V�]E�G�g��4(�y�`����?�:�S�uI��*Cy('EK����:�/�L�	�6����A���4�ǁ��o�>�ه�Эʹ:�c�W����@ A}����cݒG��%�I�(���t��I;<��i�W ��0�.��2w?��F~�h\ښb���S�ڌ3l�:<�����b�t��Jv�| e�[0`t�= ��4�0#��{x���N�Q�F�v���4҉�cӑj�gIQ*����EF��H�k"my���~h���T��]<4w�����4�(��
���5;�uD`�y�Cw��=�-�TlF�c�pm|�:�3���� ��z~���1҅E�	J%յ�b<���z:3��;2��B	G"1y?ֱ��uX�?�$l��,ʠ) �A]��
�J1T�	�v㪎�0�ة��u��AH�F�� -�*��PZ�f�_�����S���Vaje��so������f"nK"�5?����l�K�s��s]�k�/>���$���Q�ߨ���
��$�5�

��$�i�����BrNRQ��Nj��+�B���I�:5��X�N�����ܬ�B�1X	�����'��1�H�R��L$�Mf�"!<)Ua\6���a�<x]��ߘ�:�U��|���d�*z�w��t�mq!=v5�x}�ܔ��R�'J6��!A�^
 '{l]��@������g3���p|E�Y-��O��8�x�|0�fJ�ռ�A����HNׅ��LN&��w�&�{��V	�Bl�v{7�KD��%�^ aê��ëQ�`Y��P-�I�����,��JF��k������'n*�ד�ˈ���N��q�@p��;CZ���i�8�fY��(����ܗ��;dt����h���/���
N�i�gI�[�ɸqX�(:[6J����V�-���$� Y�W�FZ,d�0�{o']�@g4��V�jpQ��ezA�3�C��h`x��@�a8}�t Cu��/p	_)��������T�����+�Z{���	�<j<�ʋ�:R�ח׫(0Rh��&����}�,�O��J���1��>�0��㪑G��8��]�*^(
V��޲��$�5Q��| ��б�0�%��{`D�6u-�&��8�.��@�~��v�� 0��@�R�r��>��Ig�j��
�r��㧭ֱbۅCw��]��>�2����g��H�)��kHo{�H�Z&NBeڽb���8(�ݔW��7��"=��AF�7��o��T�n]7�~�T�i�QD��]F^D�d)�L��_`-�e��N߉����+Z�Y>QV����̻��((m���Ao��Wq�B�<0����;��[��:k#('"���7:u�wL:��a���	:���,j�,�M���V�bT�Fs����A&�Dlz�Z{󑠊6/A8Q��&u�I��]$����P ���-2ǲ�j؇��KB���ke4��]u{]Ɏ�������uU�=|U���F��s�2i��o�����&�!���h�}<{{��*���C�k��G'�M��wɽy�?����<�.�G<��|�,���!c��Dm�
�x�GD�	�i(³�H�bUz	�H��XcN��}&���7�c1*�x�f"�4��5R7�h{D;#�,p�ݑ�C����"ZV���U��?��{��DzB�AIFQ�P�EkKjP��_��d�O��p���K����ZJ���6P21��+�k���ʷx�Xئ���[���p�:\�L��g��A�:t7�"�a֕��]����XxVx����%�����a���o4`���]r��W	���iCV1Z"�]�?��+�oVza�ő\��MR�F�g��V���{ݸ��bV��rxf�G3,�)Uh���`�O��U7w)�{�<�d�m�+�.V�3��4:wFĉ��W������嚚e*Fs�m�>U�̃y�xʶٓ����tЃ׼��lF?׬�<��}��r�EjD^V�����G��qX#���&����d2�y�f��X��NB�~�����x��{�hW���xe�m��(xt��?Y���d�{�_vGPǯy����# Zܗ�z!=���WDq;"��&K���Y�F�98�mNul��k0��/ŁlKhzo&Al��w�Rؚ�<딄�3e>I����m-�sT"kiP�z��qOA�Pؽ��_D=o�Q3f��/�]��	�k�~�g��S�"��F5�
F�`mct���� ���-_*�\"�p�Lq�R����m��fe��?:�0�e4��|�^�	7�=�X�(�X/|�Sk�,sx������E�zDf�A�A�YV�������̇�_�ޔ��+ꖂcm)�96��\o*ś77daH�F�(��^�L�.���%@��~��a�x��O�G�`-�ՒH�d�$ŷaX>;m 3�|����<�@�#�'w>x�N8���ђ^4yyǉ��7F��|p��I,F<ޡˡ����؃o8�'H�iގ+d�gb~7l��pȤf\��.�����������Q��߈̬o�^j�R�����{r�npԖ+���xx��k�h"�P��!�4����D���8L>��T��S2\d�L�J�]����ޢd���8-ԜF/^`iq�,>p�+3rDtr�����t�[u�K�����C=�"F�e��.���r�}�+��Eg��n�VT̓����8�v�"e�P���+�m��ԑ�	[�<�E�_K�C�d_3����ׯ$���<��L5���W}clt��T����b�*SWCV���Kh?ǅ��	�i;u����%����B_�S�����Ӈ���T�.pF��`��r�-��,��asǨ�ܡ^ڗ�BH�=O�^'@2{�Y�4�}9�^ò+��ÞǦ@�<�O�[�nX����b�š�+�>VGy�:�	<�>i&����\��M��$���"�'}��������e�I����R����p.�y�9���=$Z�}7��2=�T��:���약���a�ӌh��y
�U���he���%�- ==�v������٪Y[��X�T�R4����h���P����p��k��o��H�����f�;�أ.&ո�~��p�ʕ(����J�J�b۞o@��]�5�B֋ �hVeؘOBI~K �p�%��u���DQ�5?#�&�2!#��,g��������1���_Ҁf-{ٯ�)�T�8.0�L�e)�Bҁ
&H��wQ�w�����@Z4��}uj�ҷ�p��:%(2�ܶ���{E��.�w����nJ�TF��Y��E1�\�A��wB����eV��
�ʄR��#WT�-j* n��
���Y��,�B�P3/8`��3��!�!.��~����=��0UI/�Uq
G�?�������o[����m(-�D�	�em¥�����Y��/�ێ�#����K�}�X�ĥ]���|�lfY΁��;ڞO�S�\�J/�n̕!��=m_���r5���ثYʢ{��m�w�i ���}x��ꨂ���Z!�k�[�j��<-cg�8M�%N���N�w����)0D3I{m����e[E�x@*)j�:��s.��@o�ǉ_��]��[h�� 1�bf���/���X���lqaD#B�?�[d������+�j{�ڡ�������nU��#�r�k��dfoqٮ������/N�=����ػ&��8�05�e��n�K�5�W�}�QU�Y��_\���9��
9U:�m8�
� *�i��"��ꗠq�]��`	h���h�E�aXL$Q�3���ǾR8B��Ж���b�-nJT~"쀔���_2`��U�_�cdE ��t�pQ�l�N,������������<ga����~�:2�\59�A����Iz�#�F-�?X�o!,�y��hs�Jm������=?g���W�3zލ��v�]p6d�7~#9ԻBu�I�v�`�����FY��K�� 	�⛼fów�Y��.�|`�wgvK�X�g�.�I�����T+^�͌�G&rsXY;�c�@s�7�'�/p���)Gg�:��@�rο���z}�_��zy�l�y�쾞�אD��r��44-;r�`�$�>��4ݧ��<m����8T��(3Ml�����տ���$2ò�9;J3rQg�`�������:��Lv�E�')f�������ԞT�;H���co�q��V�M�H���A��(�RҰ��w8�xz	�a�x�m���Ul��345[^�r�e*V4V@X%�Վ��h�t\�r���F� EE�~<9���M�b���s���Kf�w9�f����*b��	��ɴʊ �c�΃ڤ�y���t\��' [�ѝ���A~<{��Q%��3VԞ8�Lf�t�����x�dt�2�{Y����9���������rh�+|j�y�Y��Ӓ�F;{b�2� .I��R�aDèI�qy�pkl(�k��������]��@��$�A�g��$ ��5��$Id+y��D�����A��]#�Pv�jp��_"NKv���%�]�>$jq
ܸKi�Ѝ���N}�NhBJ�ȫsk��u)��b�CGdu�T���~��㤘U�KDbb�[�h�k҅��C�%גU���K��/��L�ȳ��}$��(�<�;�k��|����M�DC�E[F���0���O�˜^���؍uGj�
^�5`��Y6<�}
ź��P�h�-�  �=k���O�cv�x��5�0�jeR��B^>��� �
�`4����j������i�P'���\+�`&>����-�vd�`^���YV�D}	<�������k� �f�\\MOJ���i�ˑQQzQ�υ�g��F�t�^���ZNx�:ho��6Ϳ=T-�������+#ţo�>���b�~W�M�w/Ƣ{O����~�{&�]?��/zI~�Q4[HډT��_tyڸZM�����!o�&+9���<c����(���L�Z��*n�c�v^��ύ��w��4�}��>�z�JR�mM��s�"'��i�'�[n���m<��o��T�s�4�H�kt��Ś%�7�&༮�,�c�Z����
ze�Ij��L�{�ْ��j�Z�H��ɂ ���Y��G�����(Y(�uW�nC,sdg��N(f��LL	U6=�1�
*��(�u�+xoQ�,z�z��j���(>+Iϐߟ-s�h�n�6�ΘKt�� ��ΪiG�wp�I��~pR��Z��c�{J���0�)��
��G.�q��o�����`zԠ��ԏ�J����Z��::8��\�E���׏�y�隑��������ҷ�Lr޶�RX�b�V�~O�j���|~�����Fp����z@���e}.�R�^P�n�5����`%�~R]sǕ�.��x���*1����9E�:�A:c�Jk<�p��>(�Jj�5j�������N̩��U]T�~g�a<
9w�{tZ�*7�T�w6��Ӂk�������8���E��2(^n�/�.��\���s1��Fb6CE� cW�a
p��p�?�K
  B�0|��`�gx��Ȏ
$M�Z��S4ȃ��\+J�b�k�t�I�
��_Q^�1�%���f�"��=b�.����D;��6�J���)>>W8�d�&�5sTpV�H�a�y��֙(J�r��ӕ��d� �`��g�T�#�s�Bv��
�\�k�x���4k���؁{-�j5����C\uʐ�]R%B�"�KW��ɹt�MGa�vuyx\:���,'��ӵC+��96�Һ�(�j(�1��q��$ WԮ_vNlHa��M��2�o �7����������;yɸ�a2Wp�;�}�u���e%�0�X*\=j�(��iQ����l�ݮ�i��}3�m\�׸ϧ��,�]A��s��*� x