��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#�?�l��Z�F3~�Qp|��:��pIۄ�d�
��&��Ađĺ�M�����2�m��ahdH��I�*2L6cB��H��&�a&�sۘJ%�b��T�f�%�Kz�
�N�D�,�<!�"I��r�rJ�1M@��7ww�A��{B��Ym��ʙ�2���5>=�����Y�f�mw����Q_��!!*剘����gp�G��4�t�_Oi�q���e^9����Ok��U���bR��?��qK�d��Q2��A����uHĲ��Ks�Q�R��u ���#�S�){Y�.^+��Y�K'��r8qJ��lN82��yG�p^��lHw�� 'f\�6�G8��Gו�cc�&"�l������G��&��[MeA�a�%�tOFro�'���eW�_t/V�%�U��BȆ����$�@�z�iv�� �����wSY+D���Ʌj�f�9���gb�Qzf�/C �+�w�(���*���qQ��3�����!s.�V�߹:��{������?��� pl�Ҍe��B+v�Ӯ���l>y��X:��u@��-ܐ��ԧ�0"��"Wn?�h�FyYRXu!Ƚ����� ����Z�WԎ0� ��)��&����ҽ������p�s��iS�p�$2���7��E�G�S&� �M� 2�͘�"g�M��Q�O$�T��˾��ٿ�:z_&��eFH��|���6�׃�(m�U��[��n��=��f誨�E�Nf�i���jܙ����I$<hY��V��<SZ�o\��
�h�^��� :I�E�H�iͲ�@��0g�.-������k�/��47%eE�	�VKL�G~צ��kod�������̩�� ��*-�92u��RǤ���>#��j����[�`�#\��q����*��4��	��*���!�uؓGo���ub��n�Q�N��Q��_y��q#�kG��{	��,O,I�z�p��s@,���ϑ���H�p�ӽ(5|1�dM8���m��zl->����D���I�(�6��0�J�ۀ�,?�-`C��2J
ڞr�BE�۽t�3�B�C̉��o�#���Yb�<^h�Q�x�3A+e���_E�"P�49�Q:;���穒��F�~��14��I����OEXاl,�lf����� ��J�RF��ˎ��o���W�VAa��u\�_��x����*�ٞ�#R�A�S\��y(ڊQnx��2A�EK��#�k=�0R�4BF�gH�������:N���v'��Z�N�.EH�Wܢ�T���ﹴ�]b6>�$'�uh�;����.:J.ˇEM̙�R�i�����M��BU�[~�!�r�!��'��4K��3�y�nhP����5�w��^x��)&y�t?z��\�L�� ,�F��!m�dxX��t��#9���\�uf=N �,.;6pプ�Ò��P�ߓ���#��F�3�|6jP���'A��f��m۶�t�j�}U�]���5�������� !�A>A�:�*	@��pQ����o�����1�F呆V�G�>.�{l�Łr��+�8,����c���~�W$�\��5���)��mi�mҩid�Ù�8�+u|�X�����H��Y�~�H�!�������-0��F��1uV�SQ*V�K#�=:&��C�b��s�yc@|���r�����LBw-#@/����KiX�h�~h6��#�,���H�h��aZ����p�^7R�G5w��2�3����?g�I�f	`�.��ř���x��3�@�wm�Գ�M�����w5�u�b1�v ~��
���e��?8j�ݖm��J�'��!�k��K\Jz���JO ܈(=�����ys4o ��:����ϕ5��?9�����ul��+�O,����%��YCMXz�z��7Ǩ�6�v��A!��6*󽐳����HM���g�6$����f��X	��Д1[���إ���?����\�� "
��Hhln3�1W�Yb�z⎥}���G/���&��2�]>D����x|��ۨ�ɉd��5,N=gS&�unr5�7�=�w����"	�9��x�dIo���h�P	�t���攽R�1�lU���%F�����0�o!���ZK�t#T$����!�<0؇�9����Z�'o�^��F%g9����!�ٝ0�'N�^�>!�Fӕ�;�eps\�8��̬�7��*u4��u��i�w�RX�g��^#�Lz��C��t	�|��ab.e����b U}P�C��������*7��YB�P����dSh�߇=�K�&_q��អ/��0;�c/:�g�5�0W�1��67������W$?¥��;�F}*� 6���I��n������sf�b��2S�k!a�b�._1@K���0}!�������f��x�m�m�OFH����r"y" />լ��xq}5II�Z�����؜��SNL:����'��X����\He!�LԼ�B����'�$��Jh|���;���̺/�\��>N;���5"�� 
�X�2�j$!֓��d*����&}�Q����m��q�=j�L�D}�,���UM�_��.jr|"�غ9}�1�#mO-��_���[��^H�S?`����`���� +v)LК$SL�Y�'p_�K�ȸ��Q�R��0x%�N(zB��y/0�u�?����G�K�e����Ցh�c��z:�}�֌C��7ϒ�e��q��䍅`Yإc��&+�b���ŦM�d�9$n~�<dԥ_�c�g�)��y�5�q	WH+���kP5�a��^����Q_�|ZTu��?Lb�)�=|ޫ}���)�P;%S,��ofL_J�������n������H`������>J�K�1�ʲ���Vf��i|��q>��)�(a����]G�P�����s��Q�;�3�Q���I/YA����\��/��%n$O��)�D]�Tڄ�#�WՌ(�.ϖ:�d8�ˏt9��K4��z�{������;�C�,ɍ	gl�ԓ���,���Ѕn6���_��iea��}et��Ͻ�|���C]/�]�k�����7���:����%8�!���E��v0d M��Gj}�-31�g��2���9��KkS�����a�v��fŢ��\b㓭.�f7��]; �m_}����U��!=(m��.;e�Z�6�^:ϋ쬛ܖ��B��*g���v�I�f��,��h۹mQ��,E(�_�k#\ii8(o��f�b�K/�7	W�w*3�7Yt�N�v��*?�7d�q\k�p:ѿ١��}�#���;�P�m;��X�Ǹ���l� ��w�FDb�iA����*.�����N�]�o����ct�Nt����x� �mڪG���;��5'���a���ˉ��h�sn[E����ȃ��7��|Y^�8�S�>��Ɗ	��OHY$b����i�G��xW[�^�d=Ds��t�?��V���G힁B����")��h˅�&I�2o<�_6��J��HW4v^��*h	Q���mr�2��}�]ɉK`�G@�2���<3Bm<�c;�\�W�B�d�7��}�:^���E��B�8Rd]a�0�m3��]a��v�NP����:M��np�˨Z�%��XS��Z��D��յS��I�v�x���s��i_�oQu��f��v=*���G�B���#�۩�揜H���_�E���e"&�?*	��ŐL�����{��U��&�p!x�H��OT�ek����%E�A[ڇ]��Xm�R$��6�.���tU%m�����)d���� T�yY�0�9'4+`���N[������Sl
4ھ�v�E��Q�� co/�η�C�r`K��������s�K^����p3wh�V�Q�Gڞ��	 Ѣ~��[}|�>Ӕ��7��u�

�tT�~���okδ7������
賄�Ht�l#hM^��� "�S��뉝��9wZ��ݓ��w�,m���nk�6�[vGZ�\�foCP���Y4=Fid�V\��N��b�/,�|1��I���M�&]��H�[�`!G儔k�����	o�s+��L��䅻�v�PZz�2aI$�_�,����EA�T�+nأ&�'+�"�QM4@(�ԄC���6�1'��ql��I3��{���%Ev��2yh���r���9ڮ�B���y�9J����;>?�/|/��2@�����=YiI����]A�T(�87��[� C��H�'������'i˓��_k> ��v���t����	T�vPK�]�L��%5Λ�X!Џ9�q�f=2�4{EC�׬O�����U
��zay
Y�|6�Lp��Vņ���+���7���"�r���ʜӅ,�0�����c��%�,����Ӌ8�S��"�X�/����F�k	��s��>/����-�AÙT�H�:@�	�w���rDXY?��5 ��2���-Rta�Ʒ��*��'g��1l������):6b�[խKJ�BH�ey�V�Aj?�dQE\Z�����J�C)K��%7�Y�{�^�7{m�G7�}�F�^-��jz�<�?y���v%
�z7�.Ӈ���¥���C�����f�R�Q�6�R��=w	�˛��K�M�}]�mb;2Yx*�"����?m:��Pb�;N�e�� vz@�V
�ҁ�4~��A��''S���r=������V'~�:hߴ����b����S:�R�z��x����|�k���:�-���8��Qa����#���(�����+�o���8�p��Q�k�2+5�7�3sd���SM���ԗ�_��s�V3܁�&^p�`i��~�:��K��)��8����j�O��wUى��-�ZVa���.U��d�r���>�2�h%�Ő����0;��1���l#zs��W�_ta*��Kg�lW�&(ǻJ��� ��q,�vj��ҲZ?2��f��q��D��r2z�o�,�	��r^+EW���@E�nX��B�;w0=`�8��R6i���yӼ��/c_iǅ����}��٣�U�:�/~�+����i�ʾ���dO����s������Ǚ�S�җ��l���v����y�}=/`��Gu���?���~����
)��x��՘	�Q���o�m��eH�8=$Ai�}zc�`p{M�����N���qK�T���oF�A6w����ك�/@��!���3�
ql���u�蒏��<&TL�%�UY3�B�4��H8K�)i('EK�_��8�ZUg82�ٹT���?�e9�G���HB�鏔!�RY��e�Lq����u�Β����Z��x���N^�4�jqRN���bf�T>�9��&�p�����u�n�7	�!��˃���	��I?��z�q4�7C7��X��u���Xc�1���^�����P�>����*Ad`w��Vie�nSP�.%��OT�F�}#m�JFF�`��Ŏw���P֧�V`��	�K��2l*G�C },��ir�$yd�d����M�mͼA��FW~]gک���@0���������&���r��L�vNGW%�]���ܷ���c�F���2�ѪJ����6�1$a�|^a(�����<^'���v E#�^-ui���ѵ�S���?�vi��rL7�ǫF��7>�*>Z��w��v������R�H��c�]aߪ��Y;��@?�7U.܋;ȉ;E	ǻ��b�F0j<$=�G%��u��{jJ$��P�0c�U��U��V��ث�Öŵb��`�4 �×���}(L��zi�妏�${!�7�����H�sOi��;�ǆ�*��ߕ(��!,�o6,d�/�W��������ܡb�ɱ�ְ�t��]S/l�Q�n
����ġu�if�KE�W�0V'6�_��T,��Ȏ��%��j�yY���5��Q6��!:H�{�W�h�?V�(�l���/(:tA^J��c�5 ��+Tu%��>�/�g� 
׀�^r�|0�BY��� ����Q����;�q`�61R_
w�	���a;.�a	�HۇG�[E�[�p�UZF��@N����6���.�}3]�:M�"��(tg���{�#�״�샴�C�����ӷg��:+����;��k�3#�^���7<y{[²��E��Q0��İ��q�P������Ϳㅅ��`1��?)��Êp&5��:�d��t�kE�~9W�/��ѩ�QxK��i���d-���
��-Gh}���"CIxGWl�uJ3��ܓ��_�:>;'�܈#Z�M��ٜ#iul��}�q�w�cіE8f`Z�����
LC��DK�H�Rrs<�Q"�u0]m9�uh83�9�����m���U���[�C�)��+_u�%��R���<HS5<�����\�I>�h��*��*ů�ui���m"��-�~����+0��^v+�=��<Sc��}��!/
*?����<i���ڑ�S呠de�oF!/g!��<x�##?�0@�]�7���+��̵
�>x2�1�)x
�=�*�����(5(��O��"���r������G��캶�0�ˮc>U�n�%#�n�g�����'���
T%���1m�3v����=�H燕�^���D;+*x��sg;�0r��ZKp��&������#/�� [n"BǇ!��oA<�S�l���X^l�W����%0D��+��2w7P����"��^�f�]K��F���)�w���^I�-ȇ�gu*�ǯ�a�,��N�N��d]���7��B�;L�y&L8u���{���L�x�� ƻg]�N�$X�q�ҍ��2��f�d~�󭡑�\S���όF�}�a�9�tu���#��ٺ����f@��I��)�M��w�`��2�:=itZ0�>T,��2�b!��j����mo}����)�W�F�2a�IAe�4�]�%�� ����hEV�v�S��2�`��\vw����ёQ�a5`jg���r����@� ���&4��4(#E���|>ΐ-������duyQA�~*k���΅%������DPf\�K7L���T�� R����бK��Ӂ�(��c�nE�oe�	������%�z�`B6�NFv�P����'o9�7���8�~�O i���͉-�]��:�z��B������Oð',V$��`%��n979͟�*h�2q&˓�8����Z���!?��ҕ�qR�HM
v�ۜ\ǲ�N�ЂCl�y}ݛM��.�PZ�v����EU8����3�~RTy�	E��܁91����16����,��i��� �QO��v�Ȓ;6�but����h'�\���JJ0v�W]�ꊚL����]P�/N��b�o�l�a"N�Y~x��g4��L88�Z�8��o,c��W�k�V;Bhkl��-��6>zi��L�J��e���}�٘��ݶ��v�po���o0cA��>g���Kvu->�iB�`ujQ������wy�I���`�Z�n�vO�
r�ͺ���X
���#v�������^~�A��z�U�le/�)�
]ЅT2	�i�z5�z�1 -��*�u!A.�WQ2���FKy���������R<1�=^ +�ĆMˆ:�>�����K=�Bܑ���@���p�1C�⧺G�������/�r���u����L�C�1X����R���Gn*A1V�� W<-�K��ŗSq-\�l-MB���cA�9u}�ic�u�M�����9��n�������}s8�������<���ȕ���N}!����� ���{+!8���P���sD��T!�.�e��-�mP}^kҳy�����[�@×�"�⪚>L/��H�|�o�L�t��91��k������吔V�k�͝=�킉��Xu���<3~^W�A�]�]t�^���!�U?Z7���4j�8���OBa�{��\��{�W�.(��F��Hsme���2߁�w��*Hg����H9��+_'�����ؼ~�nv������X<�`�G���n��m�l$�������������\/.w&)��$���pf�%��̠�ŝO�?�-��L���Őo&�o�����~�Y)[���Tj��yض�*�3t���n?���Jr�:	8�^��;V^c�"������%����ݲ�!����	t˂��7C�`�0���Mh�A�Ʈ�c��-��Ll��BSbe�4�׃�Wv�H|�@e
eR���t�m�:�3�73���|�J?Au�#�����%62Z� �w�B�	����):�$<�rN���ڈ<"ݏ%���k�8+�zh(��'�4�ԉ#��?�Μ躉+ꗗ�}6�;�!IMׂ�eԁ�ퟋ{jȸ��O� ��~���u� ��H?�4��⩀�]>����z�/T�L��)Ҽ��68���i+W�[2�=��^H�6l�49�~L��M���ٰ�J�R�	��Z�٩���0r�J��֞	ɞV"�1]tT�lC�#�a`�Ĕ�R�ZPčݞ��S�\�o���a��
u'���n��z'��z�H��̙;5���,�0K}�i�̫9�MC�}iejvA&���*0��iu�W����w�}�@t��(���j�����Ƒg�Xq�D�_$��X#.͈)58�y�1����".����/�MH�1�;�ώt��q��BQ-חC���D)����UUN�?)��w�GEf`��)[�H��6���4�ZF�9W���ac�W�z��x�6r�&*I��m�9��n*~"��с؆���P�!4Ht���k��6v�ׄ,%�w��N�v��<Dx]7�;;:9����A���S"�+e�\b�{�k���E3^��K���iTt�[=ĥbp��M��Az'���9����xa�l��X^�4+�W�$�DG�
�c�ǩ��g�uG*��OM3܁z%�$�|"-�o\OJ��Ιo��c�!}�{\�l}�O=W{� ���g�J�>�z��K��`=L%�f�g@(s�"�HTĝP�5�(��'��j/)���ٽ�|j�4i�>`��/���=@q3�v~���q�WN����YQ�ɻI�f���8(�rhhU+FҺ�MK^���v�oA��)�<�)l�ֲ�3>|�.��?���"�}},l���?�W�����7�y�B)�<c�yW`RCs��C�Zߓ�Q� �r^s��1jO�[���CV�"������[H:s�ᱬ;l��=��c��ދ}��r�u�?X�~UgԵUUz�Q~d�;�𧤓��[@xF���Q,ւK"O�.	Lr\ 6|�B��S�*%6,RҼex��/'V���Z-x4H���ea�����w	�|�Z���U�G����M��Wt���k��`�a+�@��f�:�C}�������o�S&�z�`�c�:�J�C��r�Եl���H�E3��"���*�9+j�qtMB�7�Ą��t.��n#�K Zh���֒�@܇LCY�/��[e�4�4���I��#]ͧ!"�'�c�q/y#���2ނ�����9'��^㿍��'|���)8Ћ/	�U!i$��p�t"I�̩J�@��O�Y���2��63���>����4Т�b��'���s�M1-�<t�,Q4sN6&����u���OX ��TT�/~^�a���n|.D��BA)A1�Ѻ����J([jV�|w��/��5w�ď���.o����������֭��)���K�J`<4R`�3�Q�,�-M_��Kc�+>�M�S�
��)����|`�gZY�!ٚ�G&N� &��;z�;k*�`I�ڛ[w�@� 懌��V8�w�;ԫ�ƚ��_Z��S�C\@+3�7;��p��X>��U<��zڽ$�U\�3Zg�L�'+�d롫V��J�YYYi@�&��]����n����f���u=D�c��N�fϡ$���5T�-ǁ2M>�'���s�{��R�:X��hW�g�|�vOh�I�-�w4�Y��$xK�-l]��-W2+�7��c��Y�r�H*h_�U���P���K&~�\	��R���)���Y.�Sz�B�=�yj)�