��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P�|5js�[`F�q�t�(���(-jp��
�����-V�N?�;�� S���H7L���S�w�Wj�K�DP2�_K�=@�%��՜��-d֥��K��8 �R��к�u̧J�'�U,��O!`k�	vR:]L?�q�`�Oم\�y�ˆ�a燺{6����/���
�C���2�M�z1S=^�J&��7�}J���b��ĥ����g�S����j�/FY��E�ݪ��f3E/��m8������RTWq�u�AmҜNh�=P�l��"������8��mi	Jm�l5�z��&I\Y	�q��H������p�hfU���� �q3�����jG'��;���!�9�*:t�����y���o�y���Ά�_e�:�,?��nA^r#͟��x��J͋�4�g	`�o(e-�ϸ�~�f��k|�J:e�>�d�R�A�$���=�)����鶶M-�4R�QV�����Y�^���}�6�3�klI�`���	��%��/�$ü,����O�+ Q�
G�W���3�F���$�U��N�N(��j+C��$��Y�������䭺{����O�wnkg��x��G܏�7)p�>c��Aҡ���z����|�?���2ѕdp�MY�m��2��l)�^�g��`� ��=�%߉n�GdI�^5o���d��NI�.�W�i|�MD1����㖤��[@��p겍R^<%0"�Nj5��尋�G�l�q������%���j���2�y`��i��|w�3�v��ki���.������?�rg.������Rn���R�4L��zz렎�W�ɵd�3j_]�B��-�b�&��+H�F�8<@��{֮��$d%��-�UQCٰ_'8�a�r�M���:�A���"��(�_��V�x��fl�����s7��j;$7��G���#�����6N�d�����)~�\M�t4�sD�D�
�P8�\��M&OI����ᥲUT��w��s��o��p�7�p-w���R�Lӕ�ݟ�9�ss����dC]�6��o0�vޗ8��"��w���c���a�%��I��ݧl�/B\pv�Z+F�xj�2��O��܂���@�v��!�g]�0D�t��>�u���
O�v��{�Ѕo�`ӏ4Qg��f�#
v���Ʌ��0��0�$(ǂ���	�\��D�ɂ5�V�j!��k���p�D�c�5�9rUF�Rh���m]V�Ak�j�
�~�<�@���eW���fx{��rb�pF)5Ć�N�iL�<+p��v��e�O�Jq��L��Q5� d:4�a��w���M���y����Z:�
�d��&4�l|�][������]�Bw|A�!)��i��g�IS���H��+�,�%}�^m�(���{��t�0��n�>k)���Z�p��=�5��-�����:rH���2Z�!����D@�3<�fz�~J) ;oIRE~ij,�f~`_�W�Wl�]��1S�1z$���K�l��6C�ڀQ����p�Y�׏����t�ZUyl؊�XX��E��w�&�A����Ϻ�������OX�k]�kD��$��A�~(���;�����̨��+i}c>�@�8ɽ����D��j���@���6�����!2g�*��1<�,��-'
φ� V���? ώ���~�}C_ch�#f���'���~�f�Bŵ�3�u:�DH��$��J]c�:���T����X�ҷ��Ls�0}Qo4B%oI�KSo�i�X{Q�uH<�s�P�ɡ6,�Ϯ��uP�3)�v��=���lGG��f6_���R�!�v�c�t�i�d��z	H
Q|���B̄�����:i���+�ص^Uv���[�.�Z/U�t� ?O��m>	BV��z�H���%�({��\��i���:UG�xZ��h�f��r����Q#u?��iu���rC�cO�Ep�=�U���|�$W��	��hk�B$�5��Z�
�#exf�-m�g��
���@����k@jLՠu{���9Kv�c�A�P��`�4����s5���غ���3�Th��+�G}f9��>��*���y�i���b=�O� ��H�i��8Y���&R�x@���`�̳W��cO/��u{Au'/��ST�x�\p/rr0��4̦�p�O���F��Jܳ�ꅾק�?��_�t��^C��-�M;��C{hb,ƎM���k���J���){�9��M�QXq%Ȗ>�t�P|@�K�)n�u����Fʹ�Uȣ����w��F���㞬s���JWꚁ[�=�3R��N<|	i$��P�ux�m�>%��c��q�^_G����K�㰻��px2g����?�%An���b��tj�lT�Xj��kIt�U�\OhxC��D�uJ���ݱ=|3KW�啿��k \�b���2�g�<k�pX��H>K5�hWL�}_��m�7��Ǝ�	B)<Np��Tq��{4Gj�`硵���ʁ��.���y���o"���������Hj�$ՠ��%��?o-xQ�@T���P'W&���|���^B��@<�a�:1��,4���\Ս�=3�@׶�_���!C�9rݪ�2��١������Cc���!U�ySх�x/�O�V��C���m�L:��e/s��	�d�>�K���K�|�����j�߀���֔���6|5��A;�\/H��6J�k�=ţ t�ހn{�&���h{��+�Qj���aшa>�5��DQ�sp���#�nb�܇����3�n�!)�.��_��������� 5x"�;��@el#�g3�0n9�\·=���1i��QN��K���Ro�S�l'�S*v�݌b��4�I]�-��.�$6��_�E+-T��aU?B�ηed�%�кNdjk�w�).���&��^ܥ��g��'|6�QfHy7%���%�X��͸B�gF}u�.��_��0,`~�I��R�������7�uEB�Eе��Y-U��IDY3ݦK�����6���`r�� c��j[d�p8�Jfi�|����F��nrb	��L�y����\/\��t�%N�W�)|u�lv�5��<qw���I'�*�k�^܉��c���vU�������Q���d\�n'���H����%2��E�fS�z_�z�wg��EW�Vw�'�&b��R�Ppç3�����M1z-�8dȮx�:��[�$�6��v���+O��_;Yѝ��
!�>�r�R!�������Ɯ�,��"	�D�/�/ɞ��{Vq �!��7��2��CĿ-5Ef�������^׉gG�9��~ww��I��8A��Lw~�߮�*.n/F=i<S����������4�=�1s�j!�0 )������ �BVR5�N3 �CS�v�la���H8J��ȿ$�"�j9xp9����p��4�..�N�`��/8���σ)Eb落V�����(F�=Z�܍��*�Ϯ9��RBy�,��$,8B�q�[�������$8ϐZ`��B��P�ݍ+��2V}���kb8୽)^2��c��B��sd�]�֣���X�vhW��_pX:�hg���q�Noc���xٹ��H�Hɲl;��C:��K	y.f��:�*��C2@����w�#9�/�x������T��']�����;<Pn����Ӹm���%�6�5"*���������>��h�Č�,�7��uR͔�#���M�������6��ؙ�]ýF���- j,�s��%SʑR�B�O�;{'���]���I!��������D@���.6����V(r�}	����D�ؗ��T�t������۝��A��I�ŵ���bt��6F�.Qi,��0\�䮜i���Nnт��p�i>�@#��@VU����[�3�l�� m�M�v�D��:I>�*��SY�B�]QÏd���S�&mE�1h��ju�^laEg^e��ۑ����a�����pa����%�[���)Z ����bA�5L��8�E��C?����;�+����&? j-z�RIus@������N<���g^5H+��@_�/�$�n/�OAd����X_��r3�%���W����Y׳l]�*B�1��@������t��b� �n��NC؈��<]���]���xJE�q!Q�P}�ӻ;�7d�c?��s�{D��XT5�VR���M5z����gmm��������S�& ����qsr����9�=���/��s��4�ES�v��ճ���/�A�ܢ����R�4��n%��
Z�N)�)8J"p8��sa*	l��o���S�W���& _-�Fj���w@�]E+�_���2�r'�G��g��%O�-�ʟJh�^�;��Q8ڙ����n�_���AP��h�c�1����R�P�G�P��:翓Cx����a�!x��n��1݆jX��p�T��N�F�C��@�ܸ�*��G=��\�3�m���yt�Rt�*/,�}������Jz���l���]`�l۝�ơu��;�\�[s�:���A��D�֊��������ʖ�;5��%�k?�yx��ե�s����h:��uf%PT齗��K�f�"�,�M+΂y۹/�G�Q�Fu����V3�X��Y���+�r��NO��:B�k�f&v
�^���JS��Qr������Έ wC�*��0vD��Tߏ!��Y�����Q�(�4^X���}��A&��$3�W��&�-2��:�Y��kn%�y���^I+Vl�Ɓ�@k�b�A:����8���ܪ�Z-Jȇi��q��6DKA2��`*q���`~�^2�^��nQ~s������Ԟ�����=�4��R�ow�GQ$��qf}��q���������
���c�7~х����O�ŧ��՘{y>~�r(�$�+,=������~FUTq!:�ɖ��|��W<S�gmI�P	s�Z�U,��(��$Ŝ��ryd)T�e{Š��}�Y�	�*�U�;�� �c��9P���vl\�h�����憴��hB�p?��؝Yt��.�+�a���b�7ᐲ`3��Mܿύ(�ɤKNQA��!�~OX�Br�TN�mbb�T��-�y\�k9��2D��ǃ��EKO�0�ۥ�?��{���zC5����%/a�����Z�~*�֎݃"��MK�!��.0!M"vL?Xѹ���1�C�w�
L�i.��k���rj�~��f4@���k6���\N�~��� �pz~���4=UNy���d�78�_�bMgu0��:�]�2&t;�t�k){2"u�IM���ޑN��jJ�L��G΢�<Qd�e[N�΀C4*�k*�K�Yu_L����jS�����ʘ��G\J����
1>�{��ʹ8m���A�N�v������z\���L��'@�!R��=K��X�%x���X��s0
mX������DE���$�؏���=HS=yNd%{���0\Sa�������]H%8�魳�u��(�o)��W�og..[��Q�P������xz?�������3; fߏ��x�������tx�aR�,�Xj��嬜�@�=��?=�y��q�/��F�<j"��Y�6�X����,.�������(=���sR����T�@���B!���'AX�1�Lp�8�1������X�j^�68���e�[�A��;�1�.��1S&1iWw"�_
И����o��� ��{�uiaa,K{XӚ�u�A y��phO�l���$�c���(#+�@���ֽ�@y>^0��nj����\�fj�#71��>a���gy��_e��i�0,�-z���'^�F�M��X�gvt�g/VNl79]�a���.,'ɺ"`�9�_�P�٬�v�n����*����u�®7�t�>m>76��%J��`7u�K���U0��#��O�X[���W��Y��=�<<O��3,˹`t �~] i��ާ�B�&!{�w��/?�w�ܗR��w[)�p�}b��+��{O����3�L�/�:#�����u��cf��
�+5�O�G�>_N?̢<�[(��H�o(��G�ߜ�Sƻ\����e�����G%Z�g�u�Mؑ_��eUM�ސE&�	1^��ODYc�]��~��R*�����<d��Mu�� ����;��p�o4�/�Y���4��,P-�i}����9����>�'�+���n��u� ��NzV3����&Ch'�Ӗ��!�Հ=k�)n�����
R��S��/|�Q�F-�ũg�����{_��������
~���RùCRVG
�����o��[�뗫įj���g}��X����[/��{t����Hs~;�yv=+�l�ڎ��a���:�兓�e�:�h���t�B��sFy��$�]W�`�*B%��u{dH��G1^_�2&���#����R�c|���8��P,�i�I\-<���q�9�~�j�
��h��j�-`��x�@��� A�tdhY�)y���2S�3��L�zf�9xG�ŵ,�eȀt�J[JO��z�s�AhIz�>7�(��q��l���I�Ay���I�D<�_�~CI~��r��7ޢ*H_z��s߁��r$���4�@��6�9ů>Ϟ�Α2�4 [�������*��	���>!�d��C�+A�a=�5�+��ǿ�f��~!��!ѩ� �5�ek��7��3�ZC7����P�$0�7s%���9�S��ڋ�Դa����U��(�de/�
_!-�(�:��K�*宾��/damvY��~���[��#�Y2W�D_��U�g�y����}�I�sTE�F��_l5|_����( :��t��V�?%�;"�BK�<sH�{=�\��>-s��}4����J�2�yVe��-S�A.��@�eUW����e3܄��2�r�p+��M��Ϩ,�
�Έc���/�Y��\���Ͻ�-V uuj��n��nR_�1f�CC=Øifh��`���&��$C��_X��6/�E��H����D�9�g��8���@V{�# H�;��;�\W�	j87[;pٌw/G����bXݸ�����������o�5m�7H�v�W���%���J�����y�ʰzډ�-O��S��=�R�)�H�VCm�,�Z��_Ţb=�2�m�iZԥD�Ȃ�O���(�.��0�����3+�=�A&��O�R6#K2�!�`,��8�zPOr,-���=[-j,t��s��}x�s�� �Rh%�pi�<Y�l�W���4�~�%�<�g�l�^�L�ϓ��n�)���@>RU�M��!,Lp�g�y�A�y�st�ʓ-{��hS'��J��y�`���}[�r]l2�{�m����*xfH��4{�Җn�\��Y�.���ec$�x��@�s�vY�Y���x�Ij�M������v�)��U4asm\�h�V�]'މL�0{�NIuؑ��x��a�|_��Q����"|�2�i��Nj���Ad��̚����)G��R�g�$qC�<�d$�sb4O�SxbYJ�su�h�����Cƻ^&}�3��D�?��~�s	� 7mqy��ßڊZ�<����c�7�VŴ�8�۵�I� �K�@�F:�U �iZ���"%��_��&����3,X���L��5�tC��H� �YM�	Ց,��/O�Z�~��O��|�V2�d�xK��&t�D��]%z��v,\�GŹ�Q������ϔ{��}7�5d^������:tb4����A�s?�Ѕx�(�1%/=�˹���F�}�����:B۳E<y��*�˻���I_�Bb�������\Ձ�X�
�ݏ#~hb�@qm(���6x�#PnuUO�1����jխv�S��?(υ�����ȱC0��#���g|��u[gh`�J%ڥ1{5=�U����N�e�0�$`)ƨ�I�#IDԷ�}^���\	��|��y�î���]PG�*���́��b~L]W"�nI�iU$����gݥo�8Jl^��5
�&;()eH�����e(�X����r�"��]ԊF�,k�ͬƸ�WuY*���9���A��^YuM��=�㏒c;�j��~���z��30�f
�r�cs��[K��';�#�jzl��r�N{Cӌf���8�r9�����l_���E��+����Ք�:Grȡ���o�w��Jk�
�.j�v_ۧ����س?�>���<�_�;g���)Q�� ��|N������W,-�@�Z\�$��&`1y��G7y�̡���k
�M���������S�/�CN�/Q�|N�ւB`��>)��6�`�h�)6�Rشy&1�:1��?*�ґ�#�~����G/��k�C�DIL��e�5�E"�24�oc8�{j�Q�qGѥʪЌcW����=��s+.�d�/������'�p�"�z���)T��3"c���g�"��LN;]�m���+�s!���갇�$�dR;��ha�.}���j�
��>N�N�ѵ&�͜�;�~�-i�.座�3N1�v�����(�$�(w��^(ҧ�a��<T��G�A�~��4.,*�"-V$��H�&���ze�Ͻ
�3��XP�K�P1�$���o+�'��B��2F�˻���^��(��M#��^x�3~�{�eO�FU��i<y,�����qp�����U7* �>�Ͱ<=v_Wq�D�!���{��:$�!J"�l���
6?e������J:�������"�-@���:w#�
R-+����w�� =�c��#����j��Є�|@h+�{)	S�/:r�M���{���蹇��ᕽ	+T8����H�+Ó��j9�����Ƃ�Q @��Q
,	�N��O���B�@�2���!!���@�4>4Ԛz�P�&J��2Q��">e���ad����eFh.�7_9��64I89+��#�/�a�$b��|":�� =-A'�WՁ�A� �*y�|���a-���4o,���?Yk	P��MT��ߛ�-�
#S�Z� �g���Bw�U��"G��Ϛ��uX���􇳽����l���!��.h��$/�MU�j�/��L@]g�sXÓ!�pdړ1n��1�a�J��捕O�m�2��f���	��L�Խ܆_;�l���kÁ�)�w��\�K�,������y����{̕X\mv�	8<3:����� �a�Rt4ͣ�<c}d%m9�� �6��r��O�u��� ��NP�v��A����T����OL,����{��9n�c�R W����tt~Rcr����HI4��E<LB4������C���?�|�GUF3�~�f��y*�\�(��䷿b�S�,�!�& �#�d5��J��|*/����b����W�����<�3��v	�*�lB�'���L�5u9�~Av��S��
����xd[��ci`��-}�"��:�,��S�����:1�}��;)Q�f�鑽ٓx�f�j[�_��H�^�]�����U��w�DPte����l�o(�AX�/T��Ԙ>x�$�_d�V��[���h���V����O`=��4�(7�V2�+߇�KWZ���|h�a�RQM�QZ�.F���h:�u�����)-X#U�b�ޟ5!}t�֭a��o	ln�s1<�g��<�@Fp����k��ȇ:���{}|+&1r�z�,��(f�3�LG��a�;95v%D���,�V�]�����L-{����̀��o{�s�N��!��ᐠ�^6Щ(�����)��-wo _|)�!��w��0�t�<ꥃn�88�V�f�H���yUE�%��\H�S[ַD�����t�|�҄[�b���gܛ"52k*>���. r3�6)�u��ʍ�݂x� f�;��nQ����%SC3��YJ����5<�y��Q��A��Vig�3;N��ڏP��F7y87!�uQ�F0 �8b@f���=�wW�@���ڷ���O�ԓ�wm��)aUe����;�|k9���,�C�pL����6�2�y7ʛ�~յ���t�/cLrS�����.$�}���(�F�Z��GH����-�X���������\��.z3(�5m�|��%��(Z�bX���Q\L7x� �������U�W�d�i��'�<;�#2zɊ�-�^�b.�y��8^N�4U�X��\��v	_m�RBLܠda6�M���ܻ���7"6[rZ�>����|�&��.���PJ���� ��!���GP�R��.v���1�##����i�K!q*[id�yUٓ�j�`hi)��y*'dS�$��jq1����7W��$�����}��s	�B-���q~�{�D̶�3mz�z�(�3$�Q46xO0lV���=� �[ݽ�M��JƋ�;1�Ok���G�a`ǣ8q��
������Wv��N(|�d8���U.BI	�C?o.���e��������\N�SNo��7֖6ϼ�YqX.����t�y�GW
����It�$K���mXY �0�Fԧ8�\3q-�
=4���3D���#z��A�} ha�w?�IE �*d0��AuS�{�7��\O_������f4���~����
�6���妔fO�}rUu4L�]��b�� �K��Ci|z`�l�䝞�OP�e̿h� ��f΄����������_�����N�LիT�i�V�O��������Ձj���&�hճ�(B5��)k�IK~keqE.���ݭu'4�v�y�X;�T��#=�ƖR�!`��U�>������YT���d�O�ގW�g�&W��0U8-<?&v,6�N_�E65��:|�W�0�d�y��Ȳ(�Q��9f�p)������Kw���9�p���Q�c���b��/1�c�G���q���s}<����,����'v^� �S��fVTM�������ݗ�Uln2���H��n
8F��hm�OgG.�~T�_�c7��R�J����������ӫoj�qW��TV�Njr4�4'C��ʤ��oL��<��@�/:$�b+�d<{v���#��'R���/\�ZZO����g�̌��e���ԭBI������j~�qM���v�AA���tK@�����fX3a=�B1��&-�2�Ec��[&	��qtj�B����FO�QZ�1�"�3wt���Ooz��l��L�?�w��z�nx����X�$�P��y�	��M���nFU:���H�tx ��qX �m,��Q~�o���9]��:|�4G0�60�7z�7�御ȕ%��͙B���N�ޔ�-xh�N�ߌݝ,���O�.�1�-s�<��3���A�	�mΥ���v�1y������|���F�����|j�´���ɗ3�