��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P�|5js�[`F�q�t�(���(-jp��
�����-V�N?�;�� S���H7L���S�w�Wj�K�DP2�_K�=@�%��՜5�A���hD}�ϾSlI��iͮ%��h��Ԣ�^g� �lT���A�����}��LY������&�ւ#�aZ�p~�J�YGO��ra�w �_7o\���|�P�;�I8��ѣ��Y�b.'� �yh�b#�������To�{��`˄R�K)��2�Ah*��U0��<���75'��h�B�-�z�d�̮�۱�T}�?�K���ӹA���&�"�bt	]~��/���^[�;���PݴQ�$
�Z��z��&Š��s�!���
�p҈���֎&�h�
 A��Ib�D�$Q����BO	ݡC�a�L9K��ظm��s�k6�g��֭H������V�2�/��WXoI��:1K;�X�	Ǉ�`"\.#xQ9(��
U-��-��L�VS�C�P� �? ��f�?����]�YY%@�"% [G���7�pc�I�gI� g�x�y0V����`��0��IAQ.�JMqæ�1�;ߐn`���O�΋0�ticVKkY"�.:�h�.���-V�ƾ��^���R������S޾@2M}�7#~,�>l?W6Q)*#��:o�8���XS��k�
�ZQ�����9d=��I�"���Ð���ɢ��
5]���^�T��sh�tb�	����SԸ%߫�1�A�L$�h2Y2v�'��J�W��������Z[l�w}!Aέr�ʀ0]&��?$A�֐���@8����x�uB
�	('��m,� /�
G����1��=fQpW B����':��u��p-�fV��B�ƭ��*%ŸC=���b1������#ƕ�N�d���Y�60ë��_�d�� �W�������yG1�z�Q!_ֱl�04uTۮD�;�(WF!WQ�I�˅�Tf��~q�})��.�}�"��=��{7�}q��J�v��N3�Ky��0i,�:�3(-Uԍj�m�r�#��u����9�wP�Z���	ΠyGD))�	�W�ּU��wgZ�mKV4�%�^#�-� �Y"��r+o��^�ǟq���{<lج��v����i��C�\��:L�ՅI[]Q�~�(Z�c�ZM�D�� �� |ƽ6YBt�RI�С6#�D��X�rX�N��,�s�㗼n�47�;	�7���r��UrqS|����b�;�� ���^���#D��?���8Dqgd�V�z�;@�-���ެ��ͨ	Y�Xb��AO�<�WX��e��w��"�/f�8���*��q��<i��b�G=DJ�֮����`dP�y1��q'2cQ|�F"͌G�*M���&1/~2��(c���T7y����P��=J�S���f6���W��>��E��E����B��%MSA��������V����R�Ӕ*�o���n�W����}ǽ(Ԩk6�np&94溡z����U a�q��$���V.
3<MK����m��O�I�v����<?��~޸/��ӣ�g��B��٩v�9�rs "��C��Q�̋a��x�Qg� �Ϯl��T �<���+L�.+R���M����5B����f�rNB���߼�����[�.�324Z(`� �k[�g�h�]p��d�ZG9�7iq'�쫃;�؞C��R1��d��~.���ᗦ
�vx�'3�G�@L�n�8<"ׁ��,=C�dڦ��[g�U-�Rx'�(��i�6,��*J�!!��w�y��֊Wԇ���.�k�PD���Hql�\cI�}J^K)�7tgb��p���G%�@3�q��| YϿka���ő�l����8њ�=�?�؁K�V��h�@/,�����LJ�4��NE��E�x#�t�"�dq��X�q�o�qU�+�g������U�:3����h��U����W�;��% 1j1$�7�+$0�BT����5e��:։��e��@us?7���A�];d7�X���a`z�����G$8^�J\���ȴ��ɝ~����ENv����-.�q����m�W�F��W,�����3#����7�Z�j���pu�0���
��G&��u5�o2�mҁM���g;�u��'�f��B���DD��	#�4�$�Zkz��,� ����d�d�,im�0����%Ȃ2��D��=*6E'�8?��v#H@`���p���3/y]vsO�/��Ly�k�Z��>=���a��V{�D� Gg`�y�X�<Z�8�4�c/���Xt �
T��V�S�z����9c�G��x��&���Cʡ�N��m���D�#G�2�^vI�Ht���(ј˥`8G_=dW���&��Ę�������'Ķb��`�Ĉ�v|�3+�QG������H�I����/i��j&��R�K
[�K�yp1<`���o�-��cx�kCZ�;P��uT��~�Q�A�~� �wI�<�MG���v�U�ӊ����K9���s�����@R4
u8�����逎M5��!�O1~h��T���J�,`��v"_�����ο��88}+����n�Bk���_dj�����BB���/'k�r.k6my�����``���te�Qd$���8�v"��[w������Zm~��y�D�1وo�d�
o@|V�	�D��^;�(��U�t?qt�G&4,nG|�H��Z/J��dz& ��V�.H�*l����JmM�g�]q���"���?-��c�^y��{�۬����Q1Q_�����e�c1s:�ӎ�z�������S���l�OX���ZՄ�T��kM�\߱C�������up�`H<��y���|�i��Bҹ�_W2���/�Ƴ�/Z-^Y
�� 7����
q9c���W�	�Ծ1����*ztڠ����Ļb冾*�aA�Ϋ@]#�*N�'���jgo��R��W� ��b+�9� 6f#��4;A�"��v-[�	EB�S�c��3�G��5jq�Q.@?�U���[�����?a~a��ekنXgFx��"a8��@���e���p��n
^W��f�0�B����C0egI�#�O��u��m�����qXQ�S�U�z$R�N�}�{�nM���b�|�-wDQvx��^3kϺ��C*�r �
&"�W82wˑHbg񎯂 �͢P�ԉ=z���W�
4ه�c&U�mX�d�zn�̉�ͩ{-#�"�VN�:ބc�*� y��P�ͽ�sv���ɀ�uc-�}�^W9���U���r��������+�wF��2��;^�f�,C����:���b���B��1;r�uF"�/�r=����w6��t��o�K��/?UuJ��+x	Cqa���E2Ĝ���ki�Y.A��Ps؜&UЋ1�.�������H���3�#Q倢���6z��AV��1N)dժ�R��/�V˃�:F�Zx�Yτ��\T���/��Ms��jm����Mq�v���k&�I��w�X�;�\�Y�/c
 �_(���X�=��t���V�2��U�D�H��X��};|T�p'���<����x�5���հ2�O����a
5���4*���N��K��G I����q<>t��n�b�b�D��f�f%�\�Fҋ���̀E]=Qcʼ��'���~7�u�P,b؋4s;u�6��:_o�~C�]�+�$��=f���{P�l�`�ӣ�С��a������E�0�:������Ӣ������"��3�6���$�ɀt�^�I�Ϡ�����YÓ#V���h��;X3j`�J�R����?!T m�5]�p�,�<u��\���P�g�𐬴��#��7�8l��\�@P��
k'ʏR����^�<�OP1b�`��F@�u#�:Vf�v8�%NP�Q��Ǉ1�'���6��)��?�jL�C����⑯�(���}��T�'���%�}&�NB���@Tʤ!<i��*�4{2H�р4b�|�3���t�%j��6���l57.�o��x,b[�UF@���4:_F�Y��wCX{�=���)�"���Ӱg�E�YL���7.2��q��u*� VC\&c��>IV4���|�<�;���ں	�:'>�, C������@Ѳ��R�r\E���2��k	��C�V{:2�
�|BD����_9��Fr:⎁�4�kk��6�L2�ftl�Ǌ)���>�)ݲ+y�;����^���\'[�Y��^Qs�9$��lNp�~i��N��/���]�y��C��y��B+�e�R�"ݣՙ������w�.E���D�aY�%���36���k��O��N�y�u���4��qU����w�T;�3M�u��\��xP{j�t��4��7�';�X>��חA(��,o5�KN%�����Y�����Oj�/g�N'���ِ�F�U�@1��4�Ŀ���=�i*�HH���4��<�����E6Yq7R�Mʿ@���1�������:�J��Le����]j��Ze(s�M9��TD���b�!�T����	��sЮxU����o}5���]��:]L��G���g�8d��/�'i�W�Y(F/���p���r�奬��z�[��l���8z	W4{��J��l���>=Y�����ܺ�]��zHe�JD̽Իn^9)T�\�x��X�:7�������̦��*�ؿ���J�'�'����29�I�=zr�8E�#�11��i���r�E����}�A2@��\,j��rN�K���.6��~ˤ2�ܳ���o�{���L���X����6�"%�2P)t?cַ<2p�K� ���j�b������ւk�S����5*|��lC�v�T͆��q����
����A�6���׬��yXaTtCV�g��݄�^c�⽭�y󢴮ΈG�HI�Ï�Qjt@A%_��Z�
^�h����[��-���9A�1wo��F)��gl�0�^�Y�шV�ߢfYg���ǿuCs�Zm�G��gr�vJ˔��� �㩬��ӵ�h\�!Ӑ�.���K1ʔ�2�ф��.�G�\����J��:Y���Z8e/�{}� �?�N _��1��.��VmES����wB+S.���
i�B"a�qS�j֮��<F~�0:D�1j�~a��G���Z��q� �9p��`�̰-d�4j]ȫ��\���A=U�@mߓ��Τ�/R���`�>�=?BC��t������5�0D
�@W�Ұ2$���K�9�lx����p�_���`������i�mK8v��A'�Qv��$�z���*��'�Ԡzk�g����К��2��gzA��!V&4����E#�nEN7�o��p�(Q�9���)�PR;a]��֓�Q�IYV�$�b�"�<׭�)/��%g�Lu&�׶��H�!n��7�����]l�g+b���S��zSu�m���Pg��,3)���A
�t�G�S}*��!Ԥ�����$��pb����m��X^s��4f����ʕ���@��V����6�e��k�`�E������g��c�/�}�>��-���h�.�j����EHডL����OA�%�gc��0č-����-�����e�C�*�R�ƫ����~I��w����C�g�-�J u�qZ�����'�.0�3�\R��ᅨ|����
}2��>��d��7]���A���X�p\/Hèc�/ a�nL:��x˼uz��+��V�Un�	U�h�wfI"��a�]'�|-�Fg}'1�+�xYz]5v�HeCj���C�C׃��\�p�ف�M�C��l+�6n�^��I!$�&%�:�!(�_Y�eMX�2��0la�m�y��S�267z�\��W��D��I���=e�|�J{����:���N�j�53f=�M��ǭ���.�"#LO�5�Lޡ��x�WS�[=� ��!Y�Qn释�5��i$f����0Pw�]�?+��ݝ���+�n���܁�����B���y|Bi:���/��{���(��� z>dM�$4:�:Ϊ�J�� ��6A��0�c���t+�Yqc�ny�g��/��Ǩ�T��
\GRb��5�bм�؂�@��
�B�'�m�n��L+b�b���Ԭ
	ڱ;�na��A�	��"��f�X�C2��̮N|Y�%�!��B��s�h���X�1�L�[�4�c��I�]u�K��W�(B�۩UjC0H�,���"�Rӎ;T2�,�Ѩm'.�d���,�h+ F��������@^�ry"n�{��C%�����T��౩��%�@�]b45&�� y��h�Pߛ�k�_���T4�1���f�����\S��^��N��j*�NYц�8�̜S�A���R��C�y�]>����T��G���;򷾕'�5�tN��t����f7�\�>C����5��}�%��* �W�zy+gqJ��|/BV�F��EE[l��F��?�T���<;?�:s0��ʾ ih����Hf��$��A�nb$���3�yᵄN�����9ݐDQO1byo���b�L�a��@a�o �3Q%��T�v��P���>Z�ʣ�d���/X}�cŎx����e�et�[����෗��ߟo(��%N4�!N��W��={*׏�/#<ƥyX@����r��x�������mi�E�W�&X�4,ȶ���L��e�3O[����Z�X�u��|�:X�=��6��dr V$n�67�a��Cm�E3cm\�ЃCl�sdfW�n��%I�e��6t�ӚU����$��F5��_���:y��@�Fo����7&鈞,⠜�4�,EoͻIV�V/@�� H4g�o��+��v��;�aW����$���T
�}.)�7�A����ҡ���� Ǉ�����Ӂ�+Wa�m��E���޶k�jA9�j�x�|����eu��K'n@E��J���ƿw�Wq#�S3h�( �o���,��H�R�#�2N�E��Š��#�´=�&�r�7?L�DK&��-��e�S�G���p��.M�
(�ڣ�VJ$��1��L��U.���[v'�+�Mjr|/�ͥ���G������vs�����񔕸�y���U�Km]�8�3p����2�~�����6��oh0�_f����d�h	�&���CQ��p��T�;���ұr���2�)�ǣg G@�J����c+*����e	(Kg}ΪԱ���D�nŒ핤3uwv�0�u��V��׶fN�B��k���E'�Hr��-���Dx�(cD�N�����;�ؿ��q!KB�G=�Y91���^� ���"��(�:��N�m/
��@)��R����}	썌�!2\��go|bH��J���0^v�W��_���w'��| P��F�� j�!{h��J�`��
1
H����ո�o���Q�Np��y��S�l�b�a�;����ѺY��ǽ��Ip�|���%ѣbw�Y���v)m(:�C�&�d��Kǝ����iJ�)��[���ae�y�ty@�zHkRc�X��U6mW�k�����\�9���� "���q�r����E"�|-��ǒsb(�)<GO#�OIl槍��7�k�[�}z��k��I3���tO|��Z���<��+��N$UB㭗�c�%�2�J 6��|�o��o 0;����m�����Ȯ����V��lM����^�-�0��pc���� ��ő@)H�0,�gf��&9rʟD׉(����*V Y�8�f1TSF�Pߴ[a�f�iFc���C��u}3�5��M��'���$�t����:�x^�S�ء��[|�B'�<&�����3G��]�@�!��Rz!�N^��S��r�<�8��Tj k�o����UB��jY�H%�
@z�?����LRY�k�bg�>��:	��t�lK�8�İ/���{�U�� K�1���)��7����^�p����{4�����yW_/*8,/`�ˮ�t�ePR��Q�`'��d���Z�M��|׋��o@���VD/�߫^\w�����^!� ~�n6�( �п\a>oR�� ��!>����4ҷ��}?�[�$�Ģ_���'�'9������X����.����%D���(*�˷"��;�l��U�ջT���Qxs �m޵�E�����I�����q�&ɯd���M��� ��qȈ"�u�(��I)�����c��8��8N|����s���F� pN))cz[���n��(���3��FYT����]/8��:�9���a��V��*1�dJA�ɓ����dp�rD��Eh�R�þ��8���)��ܳ}�F�^�Z^��&)q�N�6@/�-Ȃ^uS����FfV�ǥ{���gnݺ</`��	�yL)n?��i��\�́F+v�s��]o
gu(��νT�
�J�K�
lW_��*�9.#����xx�gy-���7*��k�g('�>Qs4%�l&� 	Ivcmk߮����Yr	��1�2xD[�<��>}&����������
���:�.���9F֒V><1�it˺^냔]��~�\䫚�wy��`=_r #�:���`���3>��m���0?n=|zMv	q6A˶x:���~���l�`����Oc��
9���.>~��R �a}׌M1vQN�<���[s�tFK�7ꏦd�e�Y������J��s?�B4���@�C�ƣT�'Koo7�Y2Y����AƏ��7�g���� �o�&b���!1ƠNw*��51s%%��Y������L�5��,����9�+�>�{�����<3�����[O�\������_�,�w���_��T�Ce����#�J%�O�62tt�g :7��t��/��*�M�n�P�$jyå�u�%�߅�$���xW��V����q�x́�yi���?�v�@�#�|f�������U�����9N����[�U!����9[����aB/|wm<e"yt�e�^аCA�A��4J)�NkN�@"B�>�om�H 
$�=?�.��"�z���mh:RGU?*�s>iƶ��������04����Ip���Xtߒ�`�`�Gq�`E�?p*}�%8�`��(5'g�j#��C-v����0̕���\tF�b�b�yd�+u�#����aQ�Z�k�3[�5����L�o^�Ԑ1�mN�pH����:�;׬��ꭉ����\���t���_(�&C�I���%�@8G����ח/�?��ro� �`�AF�"\��ڮ���<U��2W�MmE�9C7�x���������K;�N<Gc��hu�t����)��41�/E��u��V��Q�4;�����G0Z3ڨ�Ҩ��-[�� �Ν"5	�Ge���GҠ�m��rM��8���A	4
��v����JźE`��E+��w�g�E7��_s%��gkZ���x4�몟�j��8� ��w`Vy�S�UG~�^^np�F���U蘸?���V/��4dݷ�4I��Q���`�8m�g�`h�;F+	���4�Rj�6k6��`�d�hk�������"�K>��j��H�\���ca�0���§R�����8!���T�d�˙-��yc���6�},�b"M,�"I��T�]���}4*�uX�V\��<�^`얤�T���-l�^��Ą�i�'��e ��p-��귓�<zWVlʨ��"6��KT��,`�%o��;�|<�N��5��L}G<�1V����x#���_�9Ҧb��������h ��oQq�(�(�9(\N��7�ff�9y{������deT�qR�=���"��,��S��k���Ft�]����ߙ��Y��b��%�xc���l��'����c�?,�r`�eH�ύC[��W�@gH��ʧ����iW�~�T�����x�D..B�D�l؊��d����r.,��GAZ�z,�Yk�ă����>+����s�|�y�j+���
�8 m�fQ��y?/�f~8�Yv���j���Y,����<�N OV���Ȇ�
����s\����oV�R���3{���E`��jjj�w��n�M�#�������Vw�v�o9�Q�3��pt5�`�!��A:-�CXGA��嬺���e�0.�.�����H OZϵk�������n�{��b�2
�D'(Xd�C��f.�y��ui���3ļ�&�sS�_�[��&��tH�^wZ,�s��Q�:~��r�6��۰�����ϫ"�ߠ�`�u��aVnpUtŰ��;R�2���f�h<�^tH>[䃊&�;ZF]�ϓ��}�h�5�js�V�]]��~g���vI�*�Lg�)v�O�6T@�A=�uՑ��H�^ty<b�ݘ?�Ƹ7?�b(����r
�_�nSj�����NS�J/c�J��ӄ-M�'��A&}H����1)&i��I^�R%R!�Dی���D�i������SE��K;x��ݞ	��9�۰s��cD�L��(�O�k����:~�5'�?��K�ea{"zӎ��h�I)u�4e��� �HN_2'P.%�	~��rb��Ǝ2�r]��㑃�Ա�ɞ�T-��E������s}cOF�\*�6���Fn���#0~�C�����S������m������Ws��n<��	�I"l�'����~���_{x@9![�b\�YL���,KJ]8���$8�ʯl#�2�{�J��z�0�c�O�Ĥ��kld�?�x�;Z�"XJ_��.�'+~����dP��.q9=�?�YS|�Ԉ�q}~�f�G�s�@!O��9J@����7�Ofr�ļ�������KR9��Z��[�9̄]���b(N9��̳��ϒ��{������2Ю8ѮW�9�LiYS<���_�U�4��=��B���<c��!��Z�w.�.�ΰ�7���g���>y�MVH/}����[��⟉ȝ(��7�W8�[���2Q�I�.�P��,m�����ܭ4_5GU*3����~����zT́���W�����줮k��y�ȃ�O��}��Q$$_J�_�U{sv$�b`��=J��Bl�J&Y�Knu�J�ĺ,7�h��#c2���}�`$t�aC�����6�G}�=�f2��5lw�����Im|�d�[:~�C�)���*��鎆��Btc���g����~�k+��#n��Q��H�^X|����H��d�_�ib��7Շ�Nd�K2�U���egj�y��b��K	��ĆM8�*���e�x��t��F�?!�d���-p0�<녎��F��;c�}`e{簻Z���F�j+���+�pF��V�Ü�Q�����`fbO��J5n���Yܣ�F�#]�D���(Їw��r�?k�-YVwL^�}��׊Lb>h��(Ы]�¼� �G:��4����Id��B]K�U��l��Յ�Y�[x�?� s�#g���L�'�̰$5�}1C��g��R�Õ�bg��[ Lo&�V��t˼b���3����N*7禴�4����(����O億�x氵K�G�)�@5x�8Gh�����˭M�LCz\�.�𺰫�	�6B�t��[2Zp#i��� ���F�v�p��
���=�v^��a�v���0�~d>r}P1$ί%��9�Z�7}��?�>�A!Q5�ZƯ7i$VJ�U U���0b�A���>;���G9�o!'�+�F�t���\{˖��Ѐ������F
+t�?���Ԉ��3X� p6�P����y�J6����\�+�`	X��>��s�/����o6blljjM U� ��)`�y_f�A1�(�>s�v���r����iSyq���KS|�t��$�fZ[)��Gt{�$)v�r�:!��dG�O:Q������9�k���3@\��֭���4� �L�=��⒝�pf�v��yU+�OG�3�rr|���Sx>DSS�� ��)3"�`�^��d3���/�r��.�5��J�/c�5Ǎ5�x��ZԁC�=��vJ�9��j߹,iU��1I]��_��(���߱�c���$~؈��L��,'�_���8��@���#7��D<��z�4}!%@1��4''R�k��B�]�FÖ�4B�Q�<A�n�	�}�KY���D�I	�If���3<T��+� օ9��U%P��n �c��T&y��������kFE9atн��+X���ʜ��(F�j^S�e�v��A��3�+NKHB w��Z�S�C-�P�P��]0,���k�Q�����9���;�P�f�w���2�,�q#?i�%B�h WN�Xʽ����ç
�ˈ���yR����ƼXm�Ź�>��߽���>c2���r�S�ʪ���	�F�d>B���K<�3�_�8�r�}�$�(�"���+Zm�?6
~���^�`�=��c+ �B��iN��8Iq(����wx�p�+��ឍw~wr`��1]@��~���?�6�m��!�M���X�Ѻvgy��(�tqY�A*b�P���ɦ���"*�MA� �d!o��|�p6y���3��Q�-k��k���
Fgύ�����~�h�V�MՕ��F��r�~,��z$��[5L����Y }.��w���s}�T'|�;Iz�ȹ(%!�K�����:���n�[9~�D�HP:����Y�;Ad�^������|��Ve�|Z��a������r�s�'G�l�@,~g��������Xr�g͸��G!��I��ǶF�ͣ�W9ڒ�U��t<N��6���#V+��b��m��9���d�_�`+�k�����c_��z�[[.�B�iE�Q5=A��Y�(#�ӥ��ҙ��D%�[!O�������j��C�x�����L��1����O�@����Ld�'=bV�R{A����p��u��{Z�G���[��q��窲�AجCok�Bl*
��NC#)f��b��+��e׳��Ϥ������څ��PU`m�C���~6��Ԕ.��'b:K獍���| ��4��m1O_����ѱ`�9��R�I�h|y�E�C�H�z�@���B`��D���k���(��rv�J�K�%)��?}�>]�������n�,�:K�+`�A=9������UI?�cóPT�W=�]�B_���رs>��s�$��u9�y� {#����T��j���V�S�2���~?��+v������*B�X\��bS
�`��>�b�芣};��ZԹ.�� ���S���@&t|���(��j~~��HJU��`Zo`����+��޽#�;�'0J���X��c;Y��9����+���uI�hPy�^�L���S�
� �N�rb<C�sJ��T1���(a�ܐ���W"�Ҫ`�x^PA	%XJ<���^��:g��{���!��x�:��j�ev/��ܡLI`�7C�9oz��l�i���P��_���c�~ܕ6�Q���VM�l���������&�_=r	5�m�����̇�19 �k��XcX�{-����sS��b��e����!Rv(�n;��M�o�\�7�� +!����?8��,'�H�5�3�7�C�2/��w�o�r�_C��.F7B��HU�%��C��uI̴nvv��V�R�O�������i��~b�H:��hf��w�R�3&��Ӕ�u%�F�O���`����|��)t��$?�N�>:�tek �S�p.�qG��\�Gy�mYN����|�B���&X�S^�.�Zx�O&�\mͱw*�z�5��̶�uc΋�,��]4���H�3�hx�._�֔o����r2�r����}�N���
Lo���i}	g�`�z�O>B��"2����] c���sPt���H�}����ȇZ�#��Z<�@����82
�G"�����4���+W=�l� q�0�9��Vq���zc�� ��3�e[�0�;�I���ou��V.<>�׫�'
���Zb
6�/Ì}��6h��
����W�i���D`>Կ^�˓K%9Ò0e��ȅ�:�C�TQZb˹�;��`�70H!���j�Zxy�2��Te{:b<B�)����ԅ���<�ݠ�*��-��@������_���\�+�h�
��O%'�"�f
��o��i����O���='JLf�s�/�o]��$?��
 ����M��kb�G+�!�\��\�m�e"0�YU@��|h�)&х�P ��wǏ*�4�����4ث����A��;)�Qޝ��k�]�DD�fkbL��8��f�;����KƲ�F8P\����N��r��͛q��ۨ ��柝��"D�TG�))΁#�m�;���t�گ3Od�a'��%`�T���1x�82��"�����Χs�
6��?�n�d�_IlH����\�	��<���jP�Y��KW�L�t\��JT��gP=S5&�NG��fb�徭�)A%X�8�I52��.i슟7Z,�)@�H�G�����I�\6˜�N����~Q�����="�a�Z�H1vL�ղ�)z�~��-Zՠ�As\0���;,I�zz\��c�?|���$@({�a�aqB��nc{�������j��,ߐ��F�c�T��Z��YmY���3sv�4HzhG�
j-��=*�m�wQ~/�:r9(V�k[s>�`�pI�D���� ���tw�U�EVzϋC�E�C�@����.���v�[#RY�mQ)�'�6�jp�`	�4��U��\*�ǵ�<cB��y�u�g�1�u�.��z"� �Ž����
ڞ�T�C�-�51:�n['�_㓌������Owd��!"#�7_!�O�'���+�����S��Fj�S�u�tw�%�lRǕ?&'�59,}��F�D8�	�n�7�i��V2�$3������)�"�{¶,s����U�?����w<��)��pC�	z�N�I?��A�v]���DN6��0 w��HcX<��)�q���Ӳg��x�h�d<I�����{K]��c�aE�942ua����&[h����&���u:KA{{��ZL��h��9�-W�4[|���C�F.X`Z=a>��R[̈́�C.w�&��蜊�p��9�4��U��]!;9�Ϥ����oJ��E�<�����^r���ƉnH����^ց��d�R웢6QC�ڇ`�}:��2���t�	�۽�����cUd_az�7�Ys,��;��<@!�H��(�pZ� ��lc����'CduBL]�����c�ڀ�w��ч�o�0�T�>0��6��
%+���(B�#�e��#�=��u8 7�ύ����a�.��b֕�o�e���6)!F��%:���\���q���z�%� ��T�鲡�WF��ӻT�8Z'��Jg��U*���kh��mq�g����z��o"�jwR����xOw�~��l��*T�a�������p��޷f���A7Gp@Y�D9>4��?U�z���^3=��İ�� u*����8��D�����d�V�j�]L7?��?�^D�$�}��
ׯ&���C O[�p�	y�׽h�3�p����i��kg�Bc۷3خ�6
�5����V�M10|��WrV5.?��SƯ�=�i
����}��7���j��[��܃L����{�سY�i�;����z^n��Ћ�h��[���p��Y�iF�s�ʅX����i�gl��QO
�ǁ��5͎�jyH�1f}�ݳ���?1u�r�@�8g/l�17�.�x�#!?���:�Q�y=�![�����X�il�8��O0��|7�i�2W�#��^�$��p���!�pT���/ܖ�^?���B:��l�(t%��iBt�JFf���z>�M�Z�/6�������Yq�(k��Ɖ��qr=���(7"���y������򖠳�!OZ�z��6�q��hE.�Xm`�z�����8��YgWB�g��x���'ة��w8\��1u>²���ȧ��53��+���.�tmŪ/�j�d�B�h:�N��F[��]]�
�~&��X�e_���}Y��$�K�������m��] ���EаsKJC�tۼ�C�	��40{���)(0m�~v)��^<G����M�� ��Qq\�@�[ߜ��(����7m�J 	-���C9]3Ö�-����t������_b^!�N8)Sw�y�`D�m��'��r�?�˲O{����ng;�O�M� ɋ*4 ������;�����=�K��"2c;`���d={;ŉ�a�g+j�/-�*��@���.^������c�s����[�������|�:u\B ��ZT�f5c���
Z��%	ƑY1En/������{#�"�A_��ʼ[L.$�P�~��Em)�н�_�A��r7�j�w\�d�`XţD	w��+9�-
����D���y��0|g�Ѯz_+�@�Ug=��X��;��F��2c�Z�\�i�/��S*M��h�醊7�"��fnCL��hA�T�/Xr�nn����@0����:���NL�G~P	�?	�f�h.݋��/z�#T�V5���x�C���Kj	��8���89���p2^����bS�#o��z��w��n(×җA�f��eZ�(7�I�D��A}\f^��R�Ŷ�#��D�$��L(g��n�/������-1hyҽϘ?�)�a�j��x@ͽ��oy*��+V{?e�M��0��^9�4TKQ).��"=��3��OE.�щ�Z��o�K��Z�Zt�2����@��6c�F��1������$����г�+��^��#ޭf��;�p����`�6�v@�=��oH�\����;Z:�X�9���}L%��w�'�Y��=_6�
����S�5���>`��5_;�Bn��q�$�8ش�r7s��.�do�f�3[�ʽ6����=��16]���ϋGn�'cd+���yd)�qC-2M�읎yk�{�6�o�F�i�;n~[���G:39��Tw�'zG���'Z���s��n���I~�/�����ɍH8?�^?'��7=��u���,F�SOQ3	�q2��,ǂG�GT��>R.��ww����מ����L���� �����3f~i���+X������c7�q�#�}^N�|�.0<y6�@5i���0�JxɅ
�k�T/�����[X����L�ta!47�F�9�XZu0S����l`	W�_e�4��z�\+�*�a^��B������ּu��cXes��Gg��Ⱥ\�q�`�:�Ns)��"��,8�ko����>*k.>(aD���b*��,~	����5V�"��E@<w����>�����S:��Τo:9}�.
<̝q�
c�rRj1[[R�R����J���>.a�s��#JZ���b2���T'�T�M�;�>��؍oo��~��Hʚ��3qH7#���01��r��5Ivd��- )�_�r64 d�
��%\���i@����N�ޡN�=k$��Dp
7�S;v����������oט�D^!�j�m+�/b��e�o6ܤ�q�(K|.�t1)���	�胧�JO��{��X-�0�'��PI�ӉU=���EP�t�|M�}��/��[���jS��:G\A3�6�Κ�s�w�ԏ� x q����7"�	��pP��ܐp���>�/�k#���g��{��G"�b�-l9R�8��N8�"�#���nY�P���vNO�������:F�v��3e�a$��(1�����/���5<�&��X'��q�Z���GP�L
y~щ&�����������0��Ls���P�^����<Ȏ.Z��	;�Ds�KlF}�{�_�ˊ�!���r�lC��\ǩa��Q�!	9b����3K��gQ�Nc��q;L�����Ӕ��C�Qq�	�J0��l���ݡ�R����c���>�@�b���i ����	AWil�v�l�)�;H�"뗃%j��o���0>����`PƘc�lz�E�/#*H߀W�[���N�T�Z$��D�Bg�w	]�K$Jz����N����{��>�h"�oÆ/�Y��{�"q�Qi0u\t?���5$@1�Px6������35���ް.*�� �;����?�w:Hj&h��կ��c��1x�h.���D5 oF�z(�s4�?�w��gT�D_�}����6	�c�5L0|���g��a���j��Uprm�NO�}�;�t�O��V��H	�wW��uNs�w���
�r�-��O��Z�,��z���[H�I��}-���;T7E&���&B�ᘑ�I��AF;"e�=�6W430�k]QF�$F�=$�v���7��a�)9|�je��&��Y�ex0�EI��+���WJf��B^�ǌ��!tCV-q,0SG��QiP���5���9:��M��}U���*��]nf�>F����NԀ�v�D�·bx�'�0�$��R��&�\B�?���Rh��3ka���PĐ�ܬ g	�L�S�f��P��7���ޑ�l%��\�1��r_ɿ�<j6��?1Z	��l�h�
�b���SpA�E�n]���P>)5:�i"����=�[m)5E����Ԍ	��:�M7rhz����&q�ԫΊ���"g�I#��b;ܭ �R�ru�p���j	� ���db�wV*A|<�)-<cΌP�$���~�T�Qh��4r���E��C��0�3��vÕp��^�g�{S�=k����l�]��,+F���Ōꥺ�]�����T�:p�W=6p>٨ۈ��։���8��(�Wt�ٳgq.�a�tR{V�zE�҉���K��qq����7f���H��G�9��X��c^�IW�Q���q���ɸ�YV!��$��/��&������9�f�@Eن/ʟ�-��&��b���f��~UW5�f}l�� ��IF�ؓ-ȧ��d��M����A����˱:����A2���T��W\z�*��6�^w���ٔ5�Ja��C���#�}~5�A���}��$M�uS������'N��#3�~���@
�%����-����pE�����R0���D���T� �萻�p��M����%�YqBrM�p��.t�ڴ}_��:��V�TZYa?*^!; �L�c���z����۴�c>u42�����-7�N#� %�:/+~#~��ǨH��M�?��;���ϙ0��<cXE�`��'m'�|`  6H��I�6껌��F�m�c���k��o�|(�g5�"ӨQ]�����HB�m��r{���������Ú+���?��^���^5K����@tly����-@R�*8t�z_V��r�7�[����V#>��6C�&��Ѐ��kA���{��fG��(yk�i ���3Cef�Zj}=iTH��+0���˫$�	u�;K�FA[�r��u@�-)��+���	���;}g���i3��k�w�H�t�"���=�������!���Ю P0�i�͂��x�H���94�%sZ�zb�ue���ڂ���ܬ�u砡$��r����,Ԫ}�oB��1m�������t� �$��j�A�ns�scLⳳ�״%J܁���N<w_@5K�9eł�{�:0JJB�\��G��(u����@�G�2D��SJM<��;ޓ犷9��W�6U�a�L�� U��e�{b�$�ܞ<w�EO�͎�2Ф����f�������8e�@69�x��3kl ���3+�ed�؋��]�ĸ��/�b�����-ɓ�_���B
 ���h1zw=3��?(ynw��}��M �io�1��~�&�Ù���:�5*�S
�̿�o����J�;C���Sn�D������ŭ�j%N玚:�3C�_k��k��`�.�^��5:���t\6H`Mo�Z��(��<��?���cd���*AM���1���AbZ�_���(��Ѧ����u�'�_GR���]��_urm�Ω�5.�h$�e;�M�1QI��⬲�.8��]��{v�Pw��ʧ�Bx�l�B
ƕ�&��y_
d��װv���aRFa����z�����W�
b@�c_4�Y��Y,�%��dbd��I�����٣pR�@!`b7Y�>��PyD<K�i���/t���ep� ����%�_��i��=�D�*�17	�#���^ [�R-ݫ^����Q��WX���\U�8b�Yg��
���pl��р�JH)� ��d�gԻw���ys��@���oe&�{P�Z9o�L���#������~�4���k��S��Wm����.��O��U�"'ؑdr���|�c��qԀ�(�n�Np�c��Τ*���NB��s�6�m�mm��e�c��H�9F�>��Oj�N���J��^��c��.VN���p!��,�p��1TX��fQ�	-�z}��E���R�>KS�����<����E�T~�����i��	�O���V(8����n�U�@�Jv���(
�k>p+�37�ֹ�	��������˂��"\P�^��u�e�Dp-0�<%,ܢV������P�����V�k�M� �y�g��PAJV���=�?8A�k!�P�YXn|$!d�R���4�$e�����!ʄ��U �B�HeF�59.3ډ��:4���[KC�W������2V����W�GȺ�O�*��_�n��q��������Ϟ<V)�h*�ޠK�4���&�6�������i�޼�����3_ �Wl8����C�������/ʭe�R�����]p:�|c����K��8Z�����w�	�;��HU)��4[�A�SZ���k�SB�6���'���1��E!�<��=Rs���5�J�!E\AW�`� ���O�r��HÉ��J�?���=�I�mG�b?��q��>B3��i8В�:�dܦ�G�o�� \`�d�1ux#G��o��? ˕h���r '�~a�k$;v}nh.��O�c�7���m꫁��Л��j�0��qW���e_����s^3��f��9��k�„�nw@�_5az����Lp����	`�X��qܐ<�="8��u�Q���������Լ侵��Y�2ӳ��#���qp��l�W���0eۤq����H�A�f�g�J�^�S�W�!f������7��J�~'�3V���
�0vג�}s��Y���o��z���ص�����8�6,6��QB�$7 /�c��L6�� d�Ӯ$˲�(�,p��`�������ۡR�$����=`^����>�\x�Cүs=3�3��:@QBE��d�(��ΐ)���Pw�1�SqQP�zI"�����F�b�̣�Շ+Y�.; %>!����sW�՘8|�'Z�uDs=z�P�U{��[�ӂ��g3~��ϐ�j�������3b��3���fA���}��@��/-쌱��Q��1�����1��:P����]���]�T�.^-p���S���:H����L*RW��ܡ�|p4�`���V�6����"LP�e�-�ĂLJrY� �k� ��kӉ�Kc8ލ���C9o�M<GLU�O��Ԉ����9=.+�V�yE|6��W(�ٳ��[��*<%����2�w2�Dh�?؂/��^�1���Ic���خ/��t#S�K��cF�T�E���)�HF�&�E7�b�+W?)��3�YJ�$@��:Pm|��SLZ�]���݄�����.�s�	<��DE��fX-_$���P���g�x���/��YUA6�q⢅���]��q8y����pD�1>ΣH�����[���ϙm����nLR��r�pR�(����;��ؑm0� :�i�
�ŝ]�Q�I���O�<�|2
�¾�ģ#��N�[�f�F�������m�3T�u[2U� Ƒ��߬���kA����~��|��3,\(��9ڹ}Eu��z3��]�]�-�oar��@%⣱8*�ӵ����<1�i����k��*��sJ9��͐�np��\�.Rv�VȰ�ۤ0UYQ\)�����˸���1�� ���Ǡ��`$�Ҷ+!-&p�u��υq�䩘��p�ԁ��h��CGr�B��á����]����K��J񓑀�HC'�ߣ���K�Yw����<���� �Ú�L��
��IC�����6����?��p��:9�6}�ߪ�_A������͐'~`� �h�wRG��8�CuM@eѨF�z�C�>�9<&�J,��+�ܭ{*I�Rྸ�z
ʈ�3C��e�̄0�{e������/�"����V��"��@y�����a�x�Щ�Zj�dq�7���c� H��s�Z�x�pd���
m����lsa����*:�c� săV��|�?Y��|q]���]1ݖ\!S EG��-iF���T"S�B������V;��h�V������>�Q}_+��d^��=���W$D�}r�̎�au
	 ���=4�����~55�蠲��m���@Wbwhs�q�z��|d�|V6�2�o�ʆ��|b���)�Q�� 
;��{B�����CJ�i�%���yl'O'"�}����^AN��t ��S�+䳳�"s JgY�?]�Е$�w���Y��
"���p
w�F�ptN�3��;�A�o����('³M�e-m�6�:]ĳg������(Z\�*v��J龬7+;���q�ؖ1�\;�T�$K���Y|߃���j�k�a��̭�Nmb�g|�S)t�搱�v���cҿQ6^tf86
�<�]����i��z��x��]�;�ek�G��Ly>L� �Vv��{�2r��-�½p6�D]��b�n� ��c��:M��FO���,0��&�6�ѨX<���FA牎��^V�E~� ���t���/�æ1�7��B)a�z���x�Urⷳ�v��2�����8�@J�X��(0�9` 2�׋��&=w��@a�VД��YL;��l���7�a�]��]�ϳ����]Z��U\9S0��6.�M����5�u�j��R����Bx�Ϥo�~S�����j���T��
v7bT�Nҵ���g�p	����l�i�����nO8��;���.�:"r_�<�ʹ����J��J�t}�B��鈘G>�%,�v��Wđ�`�YV�+�M����M������o�%�3��^�N�yY��|�؉y�H��5}#�4x�6��6����Q) O+Y/�^e�IW�͒u��T~��v��[����Ha\��t�T���#�=�ICb�������\c�o�(���B01"jq�/V��9QT�Gd"��� \�94���g��㞦�n[�TU�G��6�ΞVD�����T9*Z�E=,��v-�u�I�/v�$8��$ImUA,�N�wE�9u"���gܞ�'��n��&ֲXi����_1z��p�Qߙ��8y��R�k�߬��%�p�9ջ��c�Y:ҕ+�d��9@����׌iP.�J��"]�����)i��ו$9����� ��kd:EԔ�IF��Fs��A7[�ÒA�҄��:��S��6�1JËM�	KFr�l~�T�L�ޮ����zT��O�t��E��qk�7�CF:=�r6�#\�vp���"��ԜS�1�ģ:��P7��%^��QŊ���VK��J���.#�l˽e|��d�^��C(������y �=��Fx�u �C��A4���lTVŀ�g� Zy-�LF�i=���4��������sd�,�ih��#���D��s��Ht
��cӬ��:��=��|�m����@����X��S;�ѕ���HA'i4z�C�k
�Fx���r��_���Ce��g� ���'��]��t�L=�-��?�M�B�eex�{�5 �����o�U?���ё��.��I��Y�W1kq?-e1~���mC�`t���c�Fh�id/�<���(�b�Y�S��o^�;��|�R�޳�[�LBb�վe��+�Ǽ]�U��K�+<y��4����ne؟�8��G#Eұ騫,a�Y���{��A�x�Xn�.���+���zz��J��La,���j�r-�w��;1}�'Iu�RA ��@���m��y��'�U<�P�օT͇�S�ʞ�Ƃ}o&k�Rh4d̷�/K�sޠ�1�qif�y�F�$-���$V �gQN`�{
�+Xs��{Z�4�H�W�P�+�ڐ�o	j6���  .�CF����U���=V��X��C�P1�K)b��2��e�wX��Q�Jn�:�b|I�m�G����Zq��0������.z¶(���.��8������uH��bR��'�����[�R1@Q�l꾀