��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����N~@#�k�0!����+��=L���0�ԴZ�2�Mc���ZO�����=�����վ�	"cqw��a��TS[��{=:�����K��-�մ�(��k��N�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i+p���ˏ�"�`���g��!��NR�j)>���:�yP`�DSg�rd���]h&Z��^�9�a�_h���ʷ�7˿���0�_��@Ր�k�!@�(�R�P����z��{}H���_Q�hФ���]xy�0�|s��9߼L���حe=�3�����Uh=8G%�t���n�4��D�cm��zۜq�a��?w}HC�#u¨�`�L�Cަg
WS�1f�k��Z�WЁ��ehg�+ݖ��F�	Y���җ��2)W��Á$��%��-�B���C|;\�z�8����P�����`��:���\���c��E�14�QC4��l���&�d�2]JQOmF��v���'O���Q��uH��� `� ��L�Po^�6�!�p��2�er�W����,�sl7g��z4ξ^yg-<��6�,^��3�#D|�
v��P�Wz���$��C���6���p88�Hx&1>�F�+Դ�"��3��Z�	�C%<�	᪑D��_�Y�/P��Q�H�s����F	O{�o���7�sߐ(]ns�;�擺]�)�׌�e9<㨓Vo�}�7Y+B帚�G�vYO^��T
�|�����j�s@W����X�;J6W�M>#@[����<�H�����?��q�������E�	r�E&��K4��a�n��(�R(F���d�`@��Z�L��I]k��^K�?S�P���lc�q�CY��e4K$�gk��-��k&���e�²,^�+S�gaw�ҵ��(����@��an�a�4�?�-��HJ����kce��`N9��պ-E��6����-.[��eٲ���F��	5mհO?�ތ	G��K���z�:��8cU��j��1%GM9$i�ج{�+�O�h`�8�V
����ԍ��.��Dtl<��Сqs�����_�Yx�(�w�Q`�g��[�svn��H,D@6�w#�/�I+jF^͐�J�E��#|FI��'hd�xP)a��^���H��_qE��H�ϰt��^I4y�2��CKN��CT#yPHnmT�!�����B���JY ��ߦ��  �<�9���R��!����R|��q&�38�q,���VR>)B+��aE����&s�tlEy���<��ū���`�AO_Uv���ޟ�q.[{�����I��cY�G�o#,��z�.���PYh�@d�Jy��ZL[�c���M����8ġH��Ė���hUiǔ"��va?|�;�_��uJ>C�.���''�"���t�eG�i{��]�k�Bwbe`�t�#͢(�#R'�xcv�΋�C$�Z�%G�ш�][��b|ƻ~�y���&�Fcl��\?��P(q_�|�w�q�1%@X:=�V-*��Ujd�^ڳ%�i��8� FZz
��H<���Y���7]g���;��p��+!m:"C�Gv��0{�[]�-�kf��-�k+kt�ME��i�R�[��AOM*�vO�9D
I�l�ls�M>/�1uz���Sڂk�}i�c^nR�雿�?�l�̋���KE��D�G�`����@+�#J�W��_��sΤY53�_���RTJ��d+n���ø�������>CO�}p������m!ʆ[��m/@eK�.��dFǩ��~K�JT$��'��zn�H}B� }��JյƱ�u=��hEN-WEb�!K|��z���Vʯ&˦�Ю��� �b2e'	�Ǚ*<W"P�1eB�a"7���n�AHd�kN��&Sz���;3��SS��̶�km��� T��z��gk6(U���3m�e|`������"�x�X*��R����F�<�q�yk�@��U��ۅ���Eڇ���1C��	�@�����e�x���M�H��L�a� [�n^�u�Ka$e��#h��xH��n��j�-H]w'�xV��W��������gѥy��`�����b��ESV2���M��2�k��}�}��ɉז�q���tϴ�}�E@ ^팗�k���,��]���v��0�-�u3����!▕����^ i��02������������	97v/�tQᲸ�-�/b�C�q�}lZ�1^�����h���*�8�Vj�km��7Ōe��#30�{�q%�h�t(���R��to��dMQ�"2�Q�v�����ڃɎk`��y E�U��q�
��E��:�-qƲ;|:����,��l����rH�{W��h_�z���W~ta({